-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Dec 17 2017 21:46:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "timer" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of timer
entity timer is
port (
    DIGIT : out std_logic_vector(1 downto 0);
    SEG2 : out std_logic_vector(7 downto 0);
    SEG1 : out std_logic_vector(7 downto 0);
    switch_up : in std_logic;
    switch_start_stop : in std_logic;
    switch_dn : in std_logic;
    switch_cancel : in std_logic;
    CLK : in std_logic;
    BUZZER : out std_logic);
end timer;

-- Architecture of timer
-- View name is \INTERFACE\
architecture \INTERFACE\ of timer is

signal \N__14847\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \SEG1_c_5\ : std_logic;
signal \SEG1_c_6\ : std_logic;
signal \SEG1_c_4\ : std_logic;
signal \SEG1_c_3\ : std_logic;
signal \SEG1_c_1\ : std_logic;
signal \SEG1_c_2\ : std_logic;
signal \SEG1_c_0\ : std_logic;
signal \display1.prescaler8_cascade_\ : std_logic;
signal \display1.digit_dataZ0Z_3\ : std_logic;
signal \DIGIT_c_0\ : std_logic;
signal \display1.digit_dataZ0Z_2\ : std_logic;
signal \display1.digit_dataZ0Z_1\ : std_logic;
signal \display1.digit_posnZ0\ : std_logic;
signal \display1.digit_dataZ0Z_0\ : std_logic;
signal \display1.prescaler8\ : std_logic;
signal \display1.prescaler8_14\ : std_logic;
signal \display1.prescaler8_15_cascade_\ : std_logic;
signal \display1.prescaler8_21_cascade_\ : std_logic;
signal \display1.prescaler8_17_cascade_\ : std_logic;
signal \display1.prescaler8_21\ : std_logic;
signal \display1.prescaler8_17\ : std_logic;
signal \display1.prescaler8_16\ : std_logic;
signal \display1.prescaler8_13\ : std_logic;
signal \display1.prescalerZ0Z_1\ : std_logic;
signal \display1.prescalerZ0Z_0\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \display1.prescalerZ0Z_2\ : std_logic;
signal \display1.prescaler_2_cry_1\ : std_logic;
signal \display1.prescalerZ0Z_3\ : std_logic;
signal \display1.prescaler_2_cry_2\ : std_logic;
signal \display1.prescalerZ0Z_4\ : std_logic;
signal \display1.prescaler_2_4\ : std_logic;
signal \display1.prescaler_2_cry_3\ : std_logic;
signal \display1.prescalerZ0Z_5\ : std_logic;
signal \display1.prescaler_2_cry_4\ : std_logic;
signal \display1.prescalerZ0Z_6\ : std_logic;
signal \display1.prescaler_2_6\ : std_logic;
signal \display1.prescaler_2_cry_5\ : std_logic;
signal \display1.prescalerZ0Z_7\ : std_logic;
signal \display1.prescaler_2_cry_6\ : std_logic;
signal \display1.prescalerZ0Z_8\ : std_logic;
signal \display1.prescaler_2_8\ : std_logic;
signal \display1.prescaler_2_cry_7\ : std_logic;
signal \display1.prescaler_2_cry_8\ : std_logic;
signal \display1.prescalerZ0Z_9\ : std_logic;
signal \display1.prescaler_2_9\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \display1.prescaler_2_cry_9\ : std_logic;
signal \display1.prescaler_2_cry_10\ : std_logic;
signal \display1.prescaler_2_cry_11\ : std_logic;
signal \display1.prescaler_2_cry_12\ : std_logic;
signal \display1.prescalerZ0Z_14\ : std_logic;
signal \display1.prescaler_2_14\ : std_logic;
signal \display1.prescaler_2_cry_13\ : std_logic;
signal \display1.prescalerZ0Z_15\ : std_logic;
signal \display1.prescaler_2_15\ : std_logic;
signal \display1.prescaler_2_cry_14\ : std_logic;
signal \display1.prescalerZ0Z_16\ : std_logic;
signal \display1.prescaler_2_cry_15\ : std_logic;
signal \display1.prescaler_2_cry_16\ : std_logic;
signal \display1.prescalerZ0Z_17\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \display1.prescalerZ0Z_18\ : std_logic;
signal \display1.prescaler_2_cry_17\ : std_logic;
signal \display1.prescalerZ0Z_19\ : std_logic;
signal \display1.prescaler_2_cry_18\ : std_logic;
signal \display1.prescalerZ0Z_20\ : std_logic;
signal \display1.prescaler_2_cry_19\ : std_logic;
signal \display1.prescalerZ0Z_21\ : std_logic;
signal \display1.prescaler_2_cry_20\ : std_logic;
signal \display1.prescalerZ0Z_22\ : std_logic;
signal \display1.prescaler_2_cry_21\ : std_logic;
signal \display1.prescaler_2_cry_22\ : std_logic;
signal \display1.prescalerZ0Z_23\ : std_logic;
signal \display1.prescalerZ0Z_12\ : std_logic;
signal \display1.prescalerZ0Z_11\ : std_logic;
signal \display1.prescalerZ0Z_13\ : std_logic;
signal \display1.prescalerZ0Z_10\ : std_logic;
signal \display1.prescaler8_12\ : std_logic;
signal \d1.idle_i\ : std_logic;
signal \d1.trans_up_1_11_cascade_\ : std_logic;
signal \a.BUZZER3_14_cascade_\ : std_logic;
signal \a.BUZZER3_20_cascade_\ : std_logic;
signal \BUZZER_c\ : std_logic;
signal \a.BUZZER3_20\ : std_logic;
signal \a.BUZZER3_19\ : std_logic;
signal \a.BUZZER3_18\ : std_logic;
signal \a.BUZZER3_17\ : std_logic;
signal \a.BUZZER3_16_cascade_\ : std_logic;
signal \a.BUZZER3_24\ : std_logic;
signal \d1.syncZ0Z_1\ : std_logic;
signal \d1.trans_up_1_12_cascade_\ : std_logic;
signal \d1.g1_3\ : std_logic;
signal \d1.g1_4_cascade_\ : std_logic;
signal \d1.countZ0Z_1\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \d1.countZ0Z_2\ : std_logic;
signal \d1.un3_count_cry_1\ : std_logic;
signal \d1.un3_count_cry_2\ : std_logic;
signal \d1.un3_count_cry_3\ : std_logic;
signal \d1.un3_count_cry_4\ : std_logic;
signal \d1.un3_count_cry_5\ : std_logic;
signal \d1.un3_count_cry_6\ : std_logic;
signal \d1.un3_count_cry_7\ : std_logic;
signal \d1.un3_count_cry_8\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \d1.un3_count_cry_9\ : std_logic;
signal \d1.un3_count_cry_10\ : std_logic;
signal \d1.un3_count_cry_11\ : std_logic;
signal \d1.countZ0Z_13\ : std_logic;
signal \d1.un3_count_cry_12\ : std_logic;
signal \d1.countZ0Z_14\ : std_logic;
signal \d1.un3_count_cry_13\ : std_logic;
signal \d1.countZ0Z_15\ : std_logic;
signal \d1.un3_count_cry_14\ : std_logic;
signal \d1.un3_count_cry_15\ : std_logic;
signal \d1.countZ0Z_16\ : std_logic;
signal \d1.idle_i_g\ : std_logic;
signal switch_dn_c : std_logic;
signal \a.countZ0Z_1\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \a.countZ0Z_2\ : std_logic;
signal \a.count_1_cry_1\ : std_logic;
signal \a.countZ0Z_3\ : std_logic;
signal \a.count_1_cry_2\ : std_logic;
signal \a.countZ0Z_4\ : std_logic;
signal \a.count_1_cry_3\ : std_logic;
signal \a.countZ0Z_5\ : std_logic;
signal \a.count_1_cry_4\ : std_logic;
signal \a.countZ0Z_6\ : std_logic;
signal \a.count_1_cry_5\ : std_logic;
signal \a.countZ0Z_7\ : std_logic;
signal \a.count_1_cry_6\ : std_logic;
signal \a.countZ0Z_8\ : std_logic;
signal \a.count_1_8\ : std_logic;
signal \a.count_1_cry_7\ : std_logic;
signal \a.count_1_cry_8\ : std_logic;
signal \a.countZ0Z_9\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \a.countZ0Z_10\ : std_logic;
signal \a.count_1_10\ : std_logic;
signal \a.count_1_cry_9\ : std_logic;
signal \a.countZ0Z_11\ : std_logic;
signal \a.count_1_11\ : std_logic;
signal \a.count_1_cry_10\ : std_logic;
signal \a.countZ0Z_12\ : std_logic;
signal \a.count_1_12\ : std_logic;
signal \a.count_1_cry_11\ : std_logic;
signal \a.countZ0Z_13\ : std_logic;
signal \a.count_1_13\ : std_logic;
signal \a.count_1_cry_12\ : std_logic;
signal \a.countZ0Z_14\ : std_logic;
signal \a.count_1_14\ : std_logic;
signal \a.count_1_cry_13\ : std_logic;
signal \a.countZ0Z_15\ : std_logic;
signal \a.count_1_cry_14\ : std_logic;
signal \a.countZ0Z_16\ : std_logic;
signal \a.count_1_cry_15\ : std_logic;
signal \a.count_1_cry_16\ : std_logic;
signal \a.countZ0Z_17\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \a.count_1_cry_17\ : std_logic;
signal \a.count_1_cry_18\ : std_logic;
signal \a.count_1_cry_19\ : std_logic;
signal \a.count_1_cry_20\ : std_logic;
signal \a.countZ0Z_22\ : std_logic;
signal \a.count_1_cry_21\ : std_logic;
signal \a.countZ0Z_23\ : std_logic;
signal \a.count_1_cry_22\ : std_logic;
signal \a.countZ0Z_24\ : std_logic;
signal \a.count_1_cry_23\ : std_logic;
signal \a.count_1_cry_24\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \a.countZ0Z_25\ : std_logic;
signal \a.countZ0Z_18\ : std_logic;
signal \a.countZ0Z_21\ : std_logic;
signal \a.countZ0Z_20\ : std_logic;
signal \a.countZ0Z_19\ : std_logic;
signal \a.BUZZER3_15\ : std_logic;
signal \prescalerZ0Z_0\ : std_logic;
signal \prescalerZ0Z_1\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \prescalerZ0Z_2\ : std_logic;
signal prescaler_1_cry_1 : std_logic;
signal \prescalerZ0Z_3\ : std_logic;
signal prescaler_1_cry_2 : std_logic;
signal \prescalerZ0Z_4\ : std_logic;
signal prescaler_1_cry_3 : std_logic;
signal \prescalerZ0Z_5\ : std_logic;
signal prescaler_1_cry_4 : std_logic;
signal \prescalerZ0Z_6\ : std_logic;
signal prescaler_1_cry_5 : std_logic;
signal \prescalerZ0Z_7\ : std_logic;
signal prescaler_1_cry_6 : std_logic;
signal prescaler_1_cry_7 : std_logic;
signal prescaler_1_cry_8 : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal prescaler_1_cry_9 : std_logic;
signal prescaler_1_cry_10 : std_logic;
signal prescaler_1_cry_11 : std_logic;
signal prescaler_1_cry_12 : std_logic;
signal prescaler_1_cry_13 : std_logic;
signal prescaler_1_cry_14 : std_logic;
signal prescaler_1_cry_15 : std_logic;
signal prescaler_1_cry_16 : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal prescaler_1_cry_17 : std_logic;
signal prescaler_1_cry_18 : std_logic;
signal prescaler_1_cry_19 : std_logic;
signal prescaler_1_cry_20 : std_logic;
signal prescaler_1_cry_21 : std_logic;
signal prescaler_1_cry_22 : std_logic;
signal prescaler_1_cry_23 : std_logic;
signal prescaler_1_cry_24 : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal prescaler_1_cry_25 : std_logic;
signal prescaler_1_cry_26 : std_logic;
signal \prescaler_1_cry_7_THRU_CO\ : std_logic;
signal \prescalerZ0Z_8\ : std_logic;
signal \prescaler_1_cry_22_THRU_CO\ : std_logic;
signal \prescalerZ0Z_23\ : std_logic;
signal \prescaler_1_cry_23_THRU_CO\ : std_logic;
signal \prescalerZ0Z_24\ : std_logic;
signal \prescaler_1_cry_25_THRU_CO\ : std_logic;
signal \prescalerZ0Z_26\ : std_logic;
signal \prescaler_1_cry_19_THRU_CO\ : std_logic;
signal \prescaler_1_cry_20_THRU_CO\ : std_logic;
signal \prescaler_1_cry_21_THRU_CO\ : std_logic;
signal \prescaler_1_cry_12_THRU_CO\ : std_logic;
signal \prescalerZ0Z_13\ : std_logic;
signal \prescaler_1_cry_13_THRU_CO\ : std_logic;
signal \prescalerZ0Z_14\ : std_logic;
signal \prescaler_1_cry_14_THRU_CO\ : std_logic;
signal \prescalerZ0Z_15\ : std_logic;
signal \prescaler_1_cry_15_THRU_CO\ : std_logic;
signal \prescalerZ0Z_16\ : std_logic;
signal \prescaler_1_cry_17_THRU_CO\ : std_logic;
signal un1_state_3_g : std_logic;
signal \prescalerZ0Z_20\ : std_logic;
signal \prescalerZ0Z_21\ : std_logic;
signal \prescalerZ0Z_22\ : std_logic;
signal \prescalerZ0Z_18\ : std_logic;
signal decrement_time_0_prescaler10_0_and : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal decrement_time_0_prescaler10_1_and : std_logic;
signal decrement_time_0_prescaler10_0 : std_logic;
signal decrement_time_0_prescaler10_2_and : std_logic;
signal decrement_time_0_prescaler10_1 : std_logic;
signal decrement_time_0_prescaler10_3_and : std_logic;
signal decrement_time_0_prescaler10_2 : std_logic;
signal decrement_time_0_prescaler10_4_and : std_logic;
signal decrement_time_0_prescaler10_3 : std_logic;
signal decrement_time_0_prescaler10_4 : std_logic;
signal decrement_time_0_prescaler10_5 : std_logic;
signal decrement_time_0_prescaler10 : std_logic;
signal \d1.mins27_1_cascade_\ : std_logic;
signal \d1.g2Z0Z_0_cascade_\ : std_logic;
signal \d1.g0_1_a5_0_9\ : std_logic;
signal \d1.g0_1_a5_0_8\ : std_logic;
signal \d1.g0_0_0_a4_2_0\ : std_logic;
signal \d1.gZ0Z2\ : std_logic;
signal \d1.countZ0Z_0\ : std_logic;
signal \d1.countZ0Z_11\ : std_logic;
signal \d1.g2_12_0\ : std_logic;
signal \d1.g2Z0Z_12_cascade_\ : std_logic;
signal \prescalerZ0Z_10\ : std_logic;
signal \prescalerZ0Z_11\ : std_logic;
signal \prescalerZ0Z_9\ : std_logic;
signal \prescalerZ0Z_12\ : std_logic;
signal decrement_time_0_prescaler10_5_and : std_logic;
signal \prescalerZ0Z_25\ : std_logic;
signal \prescalerZ0Z_27\ : std_logic;
signal \prescalerZ0Z_17\ : std_logic;
signal \prescalerZ0Z_19\ : std_logic;
signal decrement_time_0_prescaler10_6_and : std_logic;
signal \d1.g2_7_2_cascade_\ : std_logic;
signal \d1.countZ0Z_12\ : std_logic;
signal switch_cancel_c : std_logic;
signal \d3.syncZ0Z_0\ : std_logic;
signal \d1.g2_7_1\ : std_logic;
signal \d2.syncZ0Z_0\ : std_logic;
signal \d4.idle_i\ : std_logic;
signal \d1.g2Z0Z_1_cascade_\ : std_logic;
signal \d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_\ : std_logic;
signal \a.countZ0Z_0\ : std_logic;
signal \d3.trans_up_1_15_1\ : std_logic;
signal \d3.trans_up_1_15_8\ : std_logic;
signal \d4.syncZ0Z_1\ : std_logic;
signal \d3.trans_up_1_15_7\ : std_logic;
signal \d4.trans_up_1_9\ : std_logic;
signal \d4.trans_up_1_12\ : std_logic;
signal \d4.trans_up_1_11\ : std_logic;
signal \d4.trans_up_1_13_cascade_\ : std_logic;
signal \d4.trans_up_1_10\ : std_logic;
signal \d4_trans_up_1_cascade_\ : std_logic;
signal \ten_secs_r_1_1_cascade_\ : std_logic;
signal \d3.trans_up_1_14_2_cascade_\ : std_logic;
signal \s_cancel_cascade_\ : std_logic;
signal d4_state : std_logic;
signal d4_trans_up_1 : std_logic;
signal \secs_0_sqmuxa_cascade_\ : std_logic;
signal un1_state_9_0 : std_logic;
signal \d1.ten_secs_1_sqmuxa_0\ : std_logic;
signal \d1.g2_0Z0Z_4\ : std_logic;
signal \d1.g2_0Z0Z_3\ : std_logic;
signal \ten_secs_1_sqmuxa_cascade_\ : std_logic;
signal \d1.g1_0\ : std_logic;
signal \d1.g0_0_0_0_0_cascade_\ : std_logic;
signal \mins_storedZ0Z_1\ : std_logic;
signal \d1.un1_mins_4_0_1_cascade_\ : std_logic;
signal \d1.countZ0Z_9\ : std_logic;
signal \d1.countZ0Z_8\ : std_logic;
signal \d1.countZ0Z_10\ : std_logic;
signal \d1.countZ0Z_7\ : std_logic;
signal \d1.trans_up_1_9\ : std_logic;
signal \d1.g2Z0Z_11\ : std_logic;
signal \d1.un1_mins_1_sqmuxa_0_cascade_\ : std_logic;
signal \d1.un1_mins_3_sqmuxa_0_0_cascade_\ : std_logic;
signal \d1.N_4\ : std_logic;
signal \mins_storedZ0Z_2\ : std_logic;
signal \d1.g1_cascade_\ : std_logic;
signal \d1.g1_7\ : std_logic;
signal \d1.g1_8\ : std_logic;
signal \d1.g1_14\ : std_logic;
signal \d1.g0_1_a5_0_10\ : std_logic;
signal \d1.g0_1_a5_0_15\ : std_logic;
signal \d1.trans_up_1_10\ : std_logic;
signal \d1.trans_up_1_11\ : std_logic;
signal \d1.trans_up_1_13\ : std_logic;
signal \d1.trans_up_1_0_cascade_\ : std_logic;
signal \d1.g0_2_0_o2_2_cascade_\ : std_logic;
signal \mins_storedZ0Z_0\ : std_logic;
signal \d1.g0_0_0\ : std_logic;
signal \d1.N_19_i_cascade_\ : std_logic;
signal \d1.stateZ0Z_0\ : std_logic;
signal \d1.g2_8_1\ : std_logic;
signal \d2.g0_0_10_cascade_\ : std_logic;
signal \d2.g0_0_12\ : std_logic;
signal \d2.g0_0_14_cascade_\ : std_logic;
signal \d1.g2_8_0\ : std_logic;
signal \d2.g0_0_11\ : std_logic;
signal \d2.trans_up_1_14_2\ : std_logic;
signal \d1.g2Z0Z_7_cascade_\ : std_logic;
signal \d1.g0_1_0_a4Z0Z_7_cascade_\ : std_logic;
signal \d4.countZ0Z_0\ : std_logic;
signal \d4.countZ0Z_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \d4.countZ0Z_2\ : std_logic;
signal \d4.un3_count_cry_1\ : std_logic;
signal \d4.countZ0Z_3\ : std_logic;
signal \d4.un3_count_cry_2\ : std_logic;
signal \d4.countZ0Z_4\ : std_logic;
signal \d4.un3_count_cry_3\ : std_logic;
signal \d4.countZ0Z_5\ : std_logic;
signal \d4.un3_count_cry_4\ : std_logic;
signal \d4.countZ0Z_6\ : std_logic;
signal \d4.un3_count_cry_5\ : std_logic;
signal \d4.countZ0Z_7\ : std_logic;
signal \d4.un3_count_cry_6\ : std_logic;
signal \d4.countZ0Z_8\ : std_logic;
signal \d4.un3_count_cry_7\ : std_logic;
signal \d4.un3_count_cry_8\ : std_logic;
signal \d4.countZ0Z_9\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \d4.countZ0Z_10\ : std_logic;
signal \d4.un3_count_cry_9\ : std_logic;
signal \d4.countZ0Z_11\ : std_logic;
signal \d4.un3_count_cry_10\ : std_logic;
signal \d4.countZ0Z_12\ : std_logic;
signal \d4.un3_count_cry_11\ : std_logic;
signal \d4.countZ0Z_13\ : std_logic;
signal \d4.un3_count_cry_12\ : std_logic;
signal \d4.countZ0Z_14\ : std_logic;
signal \d4.un3_count_cry_13\ : std_logic;
signal \d4.countZ0Z_15\ : std_logic;
signal \d4.un3_count_cry_14\ : std_logic;
signal \d4.un3_count_cry_15\ : std_logic;
signal \d4.countZ0Z_16\ : std_logic;
signal \d4.idle_i_g\ : std_logic;
signal \d3.countZ0Z_0\ : std_logic;
signal \d3.countZ0Z_1\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \d3.countZ0Z_2\ : std_logic;
signal \d3.un3_count_cry_1\ : std_logic;
signal \d3.countZ0Z_3\ : std_logic;
signal \d3.un3_count_cry_2\ : std_logic;
signal \d3.countZ0Z_4\ : std_logic;
signal \d3.un3_count_cry_3\ : std_logic;
signal \d3.countZ0Z_5\ : std_logic;
signal \d3.un3_count_cry_4\ : std_logic;
signal \d3.countZ0Z_6\ : std_logic;
signal \d3.un3_count_cry_5\ : std_logic;
signal \d3.countZ0Z_7\ : std_logic;
signal \d3.un3_count_cry_6\ : std_logic;
signal \d3.countZ0Z_8\ : std_logic;
signal \d3.un3_count_cry_7\ : std_logic;
signal \d3.un3_count_cry_8\ : std_logic;
signal \d3.countZ0Z_9\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \d3.countZ0Z_10\ : std_logic;
signal \d3.un3_count_cry_9\ : std_logic;
signal \d3.countZ0Z_11\ : std_logic;
signal \d3.un3_count_cry_10\ : std_logic;
signal \d3.countZ0Z_12\ : std_logic;
signal \d3.un3_count_cry_11\ : std_logic;
signal \d3.un3_count_cry_12\ : std_logic;
signal \d3.un3_count_cry_13\ : std_logic;
signal \d3.un3_count_cry_14\ : std_logic;
signal \d3.un3_count_cry_15\ : std_logic;
signal \d3.idle_i_g\ : std_logic;
signal \decrement_time_0_prescaler10_THRU_CO\ : std_logic;
signal \un1_state_7_0_cascade_\ : std_logic;
signal \un1_alarm_on_0_sqmuxa_0_i_cascade_\ : std_logic;
signal \N_120_1\ : std_logic;
signal s_cancel : std_logic;
signal \d3.countZ0Z_13\ : std_logic;
signal d3_g0_1 : std_logic;
signal \d1.secs_0_sqmuxa_xZ0Z1\ : std_logic;
signal \mins_storedZ0Z_3\ : std_logic;
signal \d1.N_5\ : std_logic;
signal \d1.un1_mins_1_sqmuxa_0\ : std_logic;
signal \d1.g0_0_0_a4_2_1\ : std_logic;
signal \secs_RNO_0Z0Z_2_cascade_\ : std_logic;
signal secs_0_sqmuxa : std_logic;
signal un1_state_7_0 : std_logic;
signal \un1_secs_c3_cascade_\ : std_logic;
signal un1_alarm_on_0_sqmuxa_0_i : std_logic;
signal \d1.trans_up_1_0\ : std_logic;
signal \d1.g2_i_a5_3\ : std_logic;
signal \d1.g0_0_0Z0Z_1_cascade_\ : std_logic;
signal \d1.g2Z0Z_10\ : std_logic;
signal \d1.g0_2_0_a4Z0Z_2\ : std_logic;
signal s_dn : std_logic;
signal \d1.g0_2_0_o2_2\ : std_logic;
signal \d1.g2_i_a5_0Z0Z_3\ : std_logic;
signal \d1.g2_i_a5_0Z0Z_6_cascade_\ : std_logic;
signal \d1.g2_i_a5Z0Z_2\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \d2.un3_count_cry_1\ : std_logic;
signal \d2.un3_count_cry_2\ : std_logic;
signal \d2.un3_count_cry_3\ : std_logic;
signal \d2.un3_count_cry_4\ : std_logic;
signal \d2.un3_count_cry_5\ : std_logic;
signal \d2.un3_count_cry_6\ : std_logic;
signal \d2.un3_count_cry_7\ : std_logic;
signal \d2.un3_count_cry_8\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \d2.un3_count_cry_9\ : std_logic;
signal \d2.un3_count_cry_10\ : std_logic;
signal \d2.un3_count_cry_11\ : std_logic;
signal \d2.un3_count_cry_12\ : std_logic;
signal \d2.un3_count_cry_13\ : std_logic;
signal \d2.un3_count_cry_14\ : std_logic;
signal \d2.un3_count_cry_15\ : std_logic;
signal \d2.idle_i_g\ : std_logic;
signal un1_state_0_sqmuxa_1_0_0 : std_logic;
signal \d1.state_1_sqmuxaZ0\ : std_logic;
signal un1_state_0_sqmuxa_1_0 : std_logic;
signal \un1_state_0_sqmuxa_1_0_cascade_\ : std_logic;
signal mins_stored_0_sqmuxa : std_logic;
signal \d1.state_0_sqmuxaZ0Z_1\ : std_logic;
signal \d1.state_0_sqmuxaZ0Z_2\ : std_logic;
signal \d1.state_0_sqmuxaZ0Z_2_cascade_\ : std_logic;
signal state_0_sqmuxa : std_logic;
signal \state_0_sqmuxa_cascade_\ : std_logic;
signal alarm_on_0_sqmuxa : std_logic;
signal \alarm_onZ0\ : std_logic;
signal \d3.countZ0Z_16\ : std_logic;
signal \d3.countZ0Z_15\ : std_logic;
signal \d3.countZ0Z_14\ : std_logic;
signal \d3.count_RNI4GDSZ0Z_16\ : std_logic;
signal \ten_secsZ0Z_2\ : std_logic;
signal un1_state_3 : std_logic;
signal \d1.g0_0Z0Z_2\ : std_logic;
signal \secsZ0Z_2\ : std_logic;
signal \secsZ0Z_1\ : std_logic;
signal \secsZ0Z_3\ : std_logic;
signal \secsZ0Z_0\ : std_logic;
signal decrement_time_0_secs9 : std_logic;
signal d2_count_6 : std_logic;
signal d2_count_5 : std_logic;
signal \d1.g2_7_0_cascade_\ : std_logic;
signal \d1.g2_11_0\ : std_logic;
signal \d1.N_3\ : std_logic;
signal \d3.trans_up_1_14_2\ : std_logic;
signal d3_trans_up_1_15 : std_logic;
signal \d1.countZ0Z_5\ : std_logic;
signal \d1.countZ0Z_4\ : std_logic;
signal \d1.countZ0Z_6\ : std_logic;
signal \d1.countZ0Z_3\ : std_logic;
signal \d1.trans_up_1_12\ : std_logic;
signal \d1.g1_9_cascade_\ : std_logic;
signal \d1.g1_13\ : std_logic;
signal un1_alarm_on_0_sqmuxa_0 : std_logic;
signal \d1.g2_iZ0Z_0\ : std_logic;
signal \d1.N_6\ : std_logic;
signal ten_secs_1_sqmuxa : std_logic;
signal \d1.mins_2_sqmuxa_1\ : std_logic;
signal \d1.mins_16_1Z0Z_3\ : std_logic;
signal \d1.g3_0_cascade_\ : std_logic;
signal \d1.N_8_0\ : std_logic;
signal mins_0_sqmuxa : std_logic;
signal \d1.g0_1_a5_0Z0Z_11\ : std_logic;
signal \d1.g2_12_1\ : std_logic;
signal d2_count_4 : std_logic;
signal d2_count_0 : std_logic;
signal \d2.trans_up_1_15\ : std_logic;
signal \d2.trans_up_1_15_cascade_\ : std_logic;
signal s_dn_0 : std_logic;
signal \d1.g2Z0Z_8\ : std_logic;
signal \d1.mins27_0_0\ : std_logic;
signal \d1.g2_i_a5_0Z0Z_7\ : std_logic;
signal d2_trans_up_1_15_1 : std_logic;
signal \d2_g0_3_cascade_\ : std_logic;
signal \d1.g2_i_a5_1Z0Z_7\ : std_logic;
signal \d2.countZ0Z_8\ : std_logic;
signal d2_trans_up_1_15_8 : std_logic;
signal \d2.countZ0Z_9\ : std_logic;
signal d2_count_16 : std_logic;
signal \d2.countZ0Z_10\ : std_logic;
signal \d2.countZ0Z_7\ : std_logic;
signal \d2.g0_0_13\ : std_logic;
signal d2_count_3 : std_logic;
signal \d1.g2_8_2\ : std_logic;
signal \d2.countZ0Z_12\ : std_logic;
signal \d2.countZ0Z_13\ : std_logic;
signal \d2.countZ0Z_14\ : std_logic;
signal \d2.countZ0Z_11\ : std_logic;
signal d2_trans_up_1_15_7 : std_logic;
signal \d1.g2_i_a5_1Z0Z_6\ : std_logic;
signal d2_sync_1 : std_logic;
signal d2_state : std_logic;
signal \d2.idle_i\ : std_logic;
signal d2_g0_3 : std_logic;
signal \d1.g0_1_0_a4Z0Z_4_cascade_\ : std_logic;
signal \stateZ0Z_1\ : std_logic;
signal \d1.g0_1_0_a4Z0Z_8\ : std_logic;
signal d2_count_15 : std_logic;
signal d2_count_2 : std_logic;
signal d2_count_1 : std_logic;
signal \stateZ0Z_0\ : std_logic;
signal \d2_g0_1_cascade_\ : std_logic;
signal \d1.g2_i_a5_1Z0Z_3\ : std_logic;
signal \d3.syncZ0Z_1\ : std_logic;
signal \d3.stateZ0\ : std_logic;
signal \d3.idle_i\ : std_logic;
signal \d1.g0_1_0Z0Z_0\ : std_logic;
signal \ten_secsZ0Z_1\ : std_logic;
signal \ten_secsZ0Z_0\ : std_logic;
signal \BNC1\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \display2.prescaler_2_cry_1\ : std_logic;
signal \display2.prescaler_2_cry_2\ : std_logic;
signal \display2.prescalerZ0Z_4\ : std_logic;
signal \display2.prescaler_2_4\ : std_logic;
signal \display2.prescaler_2_cry_3\ : std_logic;
signal \display2.prescaler_2_cry_4\ : std_logic;
signal \display2.prescalerZ0Z_6\ : std_logic;
signal \display2.prescaler_2_6\ : std_logic;
signal \display2.prescaler_2_cry_5\ : std_logic;
signal \display2.prescaler_2_cry_6\ : std_logic;
signal \display2.prescalerZ0Z_8\ : std_logic;
signal \display2.prescaler_2_8\ : std_logic;
signal \display2.prescaler_2_cry_7\ : std_logic;
signal \display2.prescaler_2_cry_8\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \display2.prescaler_2_cry_9\ : std_logic;
signal \display2.prescaler_2_cry_10\ : std_logic;
signal \display2.prescaler_2_cry_11\ : std_logic;
signal \display2.prescaler_2_cry_12\ : std_logic;
signal \display2.prescaler_2_cry_13\ : std_logic;
signal \display2.prescaler_2_cry_14\ : std_logic;
signal \display2.prescaler_2_cry_15\ : std_logic;
signal \display2.prescaler_2_cry_16\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \display2.prescaler_2_cry_17\ : std_logic;
signal \display2.prescaler_2_cry_18\ : std_logic;
signal \display2.prescaler_2_cry_19\ : std_logic;
signal \display2.prescaler_2_cry_20\ : std_logic;
signal \display2.prescaler_2_cry_21\ : std_logic;
signal \display2.prescaler_2_cry_22\ : std_logic;
signal \display2.prescalerZ0Z_23\ : std_logic;
signal \display2.prescalerZ0Z_21\ : std_logic;
signal \display2.prescalerZ0Z_20\ : std_logic;
signal \display2.prescalerZ0Z_22\ : std_logic;
signal \display2.prescalerZ0Z_19\ : std_logic;
signal \display2.prescalerZ0Z_5\ : std_logic;
signal \display2.prescalerZ0Z_3\ : std_logic;
signal \display2.prescalerZ0Z_7\ : std_logic;
signal \display2.prescalerZ0Z_2\ : std_logic;
signal \display2.prescalerZ0Z_12\ : std_logic;
signal \display2.prescalerZ0Z_10\ : std_logic;
signal \display2.prescalerZ0Z_13\ : std_logic;
signal \display2.prescalerZ0Z_11\ : std_logic;
signal \display2.prescaler8_15\ : std_logic;
signal \display2.prescaler8_12_cascade_\ : std_logic;
signal \display2.prescaler8_13\ : std_logic;
signal \display2.prescaler8_21_cascade_\ : std_logic;
signal \display2.prescalerZ0Z_1\ : std_logic;
signal \display2.prescaler8_14\ : std_logic;
signal \display2.prescaler_2_9\ : std_logic;
signal \display2.prescalerZ0Z_9\ : std_logic;
signal \display2.prescaler_2_14\ : std_logic;
signal \display2.prescalerZ0Z_14\ : std_logic;
signal \display2.prescalerZ0Z_17\ : std_logic;
signal \display2.prescalerZ0Z_16\ : std_logic;
signal \display2.prescalerZ0Z_18\ : std_logic;
signal \display2.prescalerZ0Z_0\ : std_logic;
signal \display2.prescaler8_17\ : std_logic;
signal \display2.prescaler_2_15\ : std_logic;
signal \display2.prescaler8_21\ : std_logic;
signal \display2.prescaler8_17_cascade_\ : std_logic;
signal \display2.prescaler8_16\ : std_logic;
signal \display2.prescalerZ0Z_15\ : std_logic;
signal switch_up_c : std_logic;
signal \d1.syncZ0Z_0\ : std_logic;
signal \minsZ0Z_3\ : std_logic;
signal \minsZ0Z_2\ : std_logic;
signal \minsZ0Z_1\ : std_logic;
signal \minsZ0Z_0\ : std_logic;
signal \display2.digit_posnZ0\ : std_logic;
signal \DIGIT_c_1\ : std_logic;
signal \display2.prescaler8\ : std_logic;
signal switch_start_stop_c : std_logic;
signal \d4.syncZ0Z_0\ : std_logic;
signal \SEG2_c_0\ : std_logic;
signal \SEG2_c_5\ : std_logic;
signal \SEG2_c_2\ : std_logic;
signal \SEG2_c_1\ : std_logic;
signal \SEG2_c_4\ : std_logic;
signal \SEG2_c_3\ : std_logic;
signal \display2.digit_dataZ0Z_2\ : std_logic;
signal \display2.digit_dataZ0Z_3\ : std_logic;
signal \display2.digit_dataZ0Z_1\ : std_logic;
signal \display2.digit_dataZ0Z_0\ : std_logic;
signal \SEG2_c_6\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \BUZZER_wire\ : std_logic;
signal \DIGIT_wire\ : std_logic_vector(1 downto 0);
signal \SEG1_wire\ : std_logic_vector(7 downto 0);
signal \SEG2_wire\ : std_logic_vector(7 downto 0);
signal switch_cancel_wire : std_logic;
signal switch_dn_wire : std_logic;
signal switch_start_stop_wire : std_logic;
signal switch_up_wire : std_logic;

begin
    \CLK_wire\ <= CLK;
    BUZZER <= \BUZZER_wire\;
    DIGIT <= \DIGIT_wire\;
    SEG1 <= \SEG1_wire\;
    SEG2 <= \SEG2_wire\;
    switch_cancel_wire <= switch_cancel;
    switch_dn_wire <= switch_dn;
    switch_start_stop_wire <= switch_start_stop;
    switch_up_wire <= switch_up;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__14845\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14847\,
            DIN => \N__14846\,
            DOUT => \N__14845\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14847\,
            PADOUT => \N__14846\,
            PADIN => \N__14845\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \BUZZER_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14836\,
            DIN => \N__14835\,
            DOUT => \N__14834\,
            PACKAGEPIN => \BUZZER_wire\
        );

    \BUZZER_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14836\,
            PADOUT => \N__14835\,
            PADIN => \N__14834\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6747\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DIGIT_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14827\,
            DIN => \N__14826\,
            DOUT => \N__14825\,
            PACKAGEPIN => \DIGIT_wire\(0)
        );

    \DIGIT_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14827\,
            PADOUT => \N__14826\,
            PADIN => \N__14825\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5958\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DIGIT_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14818\,
            DIN => \N__14817\,
            DOUT => \N__14816\,
            PACKAGEPIN => \DIGIT_wire\(1)
        );

    \DIGIT_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14818\,
            PADOUT => \N__14817\,
            PADIN => \N__14816\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13374\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14809\,
            DIN => \N__14808\,
            DOUT => \N__14807\,
            PACKAGEPIN => \SEG1_wire\(0)
        );

    \SEG1_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14809\,
            PADOUT => \N__14808\,
            PADIN => \N__14807\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6027\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14800\,
            DIN => \N__14799\,
            DOUT => \N__14798\,
            PACKAGEPIN => \SEG1_wire\(1)
        );

    \SEG1_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14800\,
            PADOUT => \N__14799\,
            PADIN => \N__14798\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5763\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14791\,
            DIN => \N__14790\,
            DOUT => \N__14789\,
            PACKAGEPIN => \SEG1_wire\(2)
        );

    \SEG1_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14791\,
            PADOUT => \N__14790\,
            PADIN => \N__14789\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6039\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14782\,
            DIN => \N__14781\,
            DOUT => \N__14780\,
            PACKAGEPIN => \SEG1_wire\(3)
        );

    \SEG1_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14782\,
            PADOUT => \N__14781\,
            PADIN => \N__14780\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5772\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14773\,
            DIN => \N__14772\,
            DOUT => \N__14771\,
            PACKAGEPIN => \SEG1_wire\(4)
        );

    \SEG1_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14773\,
            PADOUT => \N__14772\,
            PADIN => \N__14771\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5781\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14764\,
            DIN => \N__14763\,
            DOUT => \N__14762\,
            PACKAGEPIN => \SEG1_wire\(5)
        );

    \SEG1_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14764\,
            PADOUT => \N__14763\,
            PADIN => \N__14762\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5811\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14755\,
            DIN => \N__14754\,
            DOUT => \N__14753\,
            PACKAGEPIN => \SEG1_wire\(6)
        );

    \SEG1_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14755\,
            PADOUT => \N__14754\,
            PADIN => \N__14753\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5796\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG1_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14746\,
            DIN => \N__14745\,
            DOUT => \N__14744\,
            PACKAGEPIN => \SEG1_wire\(7)
        );

    \SEG1_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14746\,
            PADOUT => \N__14745\,
            PADIN => \N__14744\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14737\,
            DIN => \N__14736\,
            DOUT => \N__14735\,
            PACKAGEPIN => \SEG2_wire\(0)
        );

    \SEG2_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14737\,
            PADOUT => \N__14736\,
            PADIN => \N__14735\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13299\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14728\,
            DIN => \N__14727\,
            DOUT => \N__14726\,
            PACKAGEPIN => \SEG2_wire\(1)
        );

    \SEG2_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14728\,
            PADOUT => \N__14727\,
            PADIN => \N__14726\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14589\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14719\,
            DIN => \N__14718\,
            DOUT => \N__14717\,
            PACKAGEPIN => \SEG2_wire\(2)
        );

    \SEG2_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14719\,
            PADOUT => \N__14718\,
            PADIN => \N__14717\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14601\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14710\,
            DIN => \N__14709\,
            DOUT => \N__14708\,
            PACKAGEPIN => \SEG2_wire\(3)
        );

    \SEG2_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14710\,
            PADOUT => \N__14709\,
            PADIN => \N__14708\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14559\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14701\,
            DIN => \N__14700\,
            DOUT => \N__14699\,
            PACKAGEPIN => \SEG2_wire\(4)
        );

    \SEG2_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14701\,
            PADOUT => \N__14700\,
            PADIN => \N__14699\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14574\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14692\,
            DIN => \N__14691\,
            DOUT => \N__14690\,
            PACKAGEPIN => \SEG2_wire\(5)
        );

    \SEG2_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14692\,
            PADOUT => \N__14691\,
            PADIN => \N__14690\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14619\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14683\,
            DIN => \N__14682\,
            DOUT => \N__14681\,
            PACKAGEPIN => \SEG2_wire\(6)
        );

    \SEG2_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14683\,
            PADOUT => \N__14682\,
            PADIN => \N__14681\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14295\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \SEG2_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14674\,
            DIN => \N__14673\,
            DOUT => \N__14672\,
            PACKAGEPIN => \SEG2_wire\(7)
        );

    \SEG2_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14674\,
            PADOUT => \N__14673\,
            PADIN => \N__14672\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_cancel_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14665\,
            DIN => \N__14664\,
            DOUT => \N__14663\,
            PACKAGEPIN => switch_cancel_wire
        );

    \switch_cancel_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14665\,
            PADOUT => \N__14664\,
            PADIN => \N__14663\,
            CLOCKENABLE => 'H',
            DIN0 => switch_cancel_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_dn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14656\,
            DIN => \N__14655\,
            DOUT => \N__14654\,
            PACKAGEPIN => switch_dn_wire
        );

    \switch_dn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14656\,
            PADOUT => \N__14655\,
            PADIN => \N__14654\,
            CLOCKENABLE => 'H',
            DIN0 => switch_dn_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14647\,
            DIN => \N__14646\,
            DOUT => \N__14645\,
            PACKAGEPIN => switch_start_stop_wire
        );

    \switch_start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14647\,
            PADOUT => \N__14646\,
            PADIN => \N__14645\,
            CLOCKENABLE => 'H',
            DIN0 => switch_start_stop_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_up_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14638\,
            DIN => \N__14637\,
            DOUT => \N__14636\,
            PACKAGEPIN => switch_up_wire
        );

    \switch_up_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14638\,
            PADOUT => \N__14637\,
            PADIN => \N__14636\,
            CLOCKENABLE => 'H',
            DIN0 => switch_up_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__3446\ : IoInMux
    port map (
            O => \N__14619\,
            I => \N__14616\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__14616\,
            I => \N__14613\
        );

    \I__3444\ : Span4Mux_s2_h
    port map (
            O => \N__14613\,
            I => \N__14610\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__14610\,
            I => \N__14607\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__14607\,
            I => \N__14604\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__14604\,
            I => \SEG2_c_5\
        );

    \I__3440\ : IoInMux
    port map (
            O => \N__14601\,
            I => \N__14598\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__14598\,
            I => \N__14595\
        );

    \I__3438\ : Span4Mux_s3_h
    port map (
            O => \N__14595\,
            I => \N__14592\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__14592\,
            I => \SEG2_c_2\
        );

    \I__3436\ : IoInMux
    port map (
            O => \N__14589\,
            I => \N__14586\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__14586\,
            I => \N__14583\
        );

    \I__3434\ : IoSpan4Mux
    port map (
            O => \N__14583\,
            I => \N__14580\
        );

    \I__3433\ : Span4Mux_s3_h
    port map (
            O => \N__14580\,
            I => \N__14577\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__14577\,
            I => \SEG2_c_1\
        );

    \I__3431\ : IoInMux
    port map (
            O => \N__14574\,
            I => \N__14571\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__14571\,
            I => \N__14568\
        );

    \I__3429\ : IoSpan4Mux
    port map (
            O => \N__14568\,
            I => \N__14565\
        );

    \I__3428\ : Span4Mux_s2_h
    port map (
            O => \N__14565\,
            I => \N__14562\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__14562\,
            I => \SEG2_c_4\
        );

    \I__3426\ : IoInMux
    port map (
            O => \N__14559\,
            I => \N__14556\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__3424\ : IoSpan4Mux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__3423\ : Span4Mux_s3_h
    port map (
            O => \N__14550\,
            I => \N__14547\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__14547\,
            I => \SEG2_c_3\
        );

    \I__3421\ : InMux
    port map (
            O => \N__14544\,
            I => \N__14534\
        );

    \I__3420\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14534\
        );

    \I__3419\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14534\
        );

    \I__3418\ : InMux
    port map (
            O => \N__14541\,
            I => \N__14531\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__14534\,
            I => \N__14528\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__14531\,
            I => \N__14525\
        );

    \I__3415\ : Span4Mux_h
    port map (
            O => \N__14528\,
            I => \N__14518\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__14525\,
            I => \N__14515\
        );

    \I__3413\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14510\
        );

    \I__3412\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14510\
        );

    \I__3411\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14507\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__14521\,
            I => \N__14504\
        );

    \I__3409\ : Span4Mux_h
    port map (
            O => \N__14518\,
            I => \N__14501\
        );

    \I__3408\ : Sp12to4
    port map (
            O => \N__14515\,
            I => \N__14494\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__14510\,
            I => \N__14494\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__14507\,
            I => \N__14494\
        );

    \I__3405\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14491\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__14501\,
            I => \display2.digit_dataZ0Z_2\
        );

    \I__3403\ : Odrv12
    port map (
            O => \N__14494\,
            I => \display2.digit_dataZ0Z_2\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__14491\,
            I => \display2.digit_dataZ0Z_2\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__14484\,
            I => \N__14481\
        );

    \I__3400\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14469\
        );

    \I__3399\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14469\
        );

    \I__3398\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14469\
        );

    \I__3397\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14466\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__14477\,
            I => \N__14462\
        );

    \I__3395\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14458\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__14469\,
            I => \N__14453\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__14466\,
            I => \N__14453\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14450\
        );

    \I__3391\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14445\
        );

    \I__3390\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14445\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__14458\,
            I => \N__14440\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__14453\,
            I => \N__14440\
        );

    \I__3387\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14437\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__14445\,
            I => \N__14434\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__14440\,
            I => \N__14431\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__14437\,
            I => \display2.digit_dataZ0Z_3\
        );

    \I__3383\ : Odrv12
    port map (
            O => \N__14434\,
            I => \display2.digit_dataZ0Z_3\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__14431\,
            I => \display2.digit_dataZ0Z_3\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__14424\,
            I => \N__14419\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__14423\,
            I => \N__14416\
        );

    \I__3379\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14411\
        );

    \I__3378\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14411\
        );

    \I__3377\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14408\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__14411\,
            I => \N__14402\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14399\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__14407\,
            I => \N__14396\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__14406\,
            I => \N__14392\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__14405\,
            I => \N__14389\
        );

    \I__3371\ : Span4Mux_v
    port map (
            O => \N__14402\,
            I => \N__14385\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__14399\,
            I => \N__14382\
        );

    \I__3369\ : InMux
    port map (
            O => \N__14396\,
            I => \N__14375\
        );

    \I__3368\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14375\
        );

    \I__3367\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14375\
        );

    \I__3366\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14372\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__14388\,
            I => \N__14369\
        );

    \I__3364\ : Sp12to4
    port map (
            O => \N__14385\,
            I => \N__14360\
        );

    \I__3363\ : Sp12to4
    port map (
            O => \N__14382\,
            I => \N__14360\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__14375\,
            I => \N__14360\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__14372\,
            I => \N__14360\
        );

    \I__3360\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14357\
        );

    \I__3359\ : Odrv12
    port map (
            O => \N__14360\,
            I => \display2.digit_dataZ0Z_1\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__14357\,
            I => \display2.digit_dataZ0Z_1\
        );

    \I__3357\ : InMux
    port map (
            O => \N__14352\,
            I => \N__14345\
        );

    \I__3356\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14345\
        );

    \I__3355\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14342\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__14345\,
            I => \N__14339\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14336\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14328\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__14336\,
            I => \N__14325\
        );

    \I__3350\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14318\
        );

    \I__3349\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14318\
        );

    \I__3348\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14318\
        );

    \I__3347\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14315\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__14331\,
            I => \N__14312\
        );

    \I__3345\ : Sp12to4
    port map (
            O => \N__14328\,
            I => \N__14303\
        );

    \I__3344\ : Sp12to4
    port map (
            O => \N__14325\,
            I => \N__14303\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__14318\,
            I => \N__14303\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__14315\,
            I => \N__14303\
        );

    \I__3341\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14300\
        );

    \I__3340\ : Odrv12
    port map (
            O => \N__14303\,
            I => \display2.digit_dataZ0Z_0\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__14300\,
            I => \display2.digit_dataZ0Z_0\
        );

    \I__3338\ : IoInMux
    port map (
            O => \N__14295\,
            I => \N__14292\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__14292\,
            I => \N__14289\
        );

    \I__3336\ : Span4Mux_s3_h
    port map (
            O => \N__14289\,
            I => \N__14286\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__14286\,
            I => \N__14283\
        );

    \I__3334\ : Span4Mux_v
    port map (
            O => \N__14283\,
            I => \N__14280\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__14280\,
            I => \SEG2_c_6\
        );

    \I__3332\ : ClkMux
    port map (
            O => \N__14277\,
            I => \N__14055\
        );

    \I__3331\ : ClkMux
    port map (
            O => \N__14276\,
            I => \N__14055\
        );

    \I__3330\ : ClkMux
    port map (
            O => \N__14275\,
            I => \N__14055\
        );

    \I__3329\ : ClkMux
    port map (
            O => \N__14274\,
            I => \N__14055\
        );

    \I__3328\ : ClkMux
    port map (
            O => \N__14273\,
            I => \N__14055\
        );

    \I__3327\ : ClkMux
    port map (
            O => \N__14272\,
            I => \N__14055\
        );

    \I__3326\ : ClkMux
    port map (
            O => \N__14271\,
            I => \N__14055\
        );

    \I__3325\ : ClkMux
    port map (
            O => \N__14270\,
            I => \N__14055\
        );

    \I__3324\ : ClkMux
    port map (
            O => \N__14269\,
            I => \N__14055\
        );

    \I__3323\ : ClkMux
    port map (
            O => \N__14268\,
            I => \N__14055\
        );

    \I__3322\ : ClkMux
    port map (
            O => \N__14267\,
            I => \N__14055\
        );

    \I__3321\ : ClkMux
    port map (
            O => \N__14266\,
            I => \N__14055\
        );

    \I__3320\ : ClkMux
    port map (
            O => \N__14265\,
            I => \N__14055\
        );

    \I__3319\ : ClkMux
    port map (
            O => \N__14264\,
            I => \N__14055\
        );

    \I__3318\ : ClkMux
    port map (
            O => \N__14263\,
            I => \N__14055\
        );

    \I__3317\ : ClkMux
    port map (
            O => \N__14262\,
            I => \N__14055\
        );

    \I__3316\ : ClkMux
    port map (
            O => \N__14261\,
            I => \N__14055\
        );

    \I__3315\ : ClkMux
    port map (
            O => \N__14260\,
            I => \N__14055\
        );

    \I__3314\ : ClkMux
    port map (
            O => \N__14259\,
            I => \N__14055\
        );

    \I__3313\ : ClkMux
    port map (
            O => \N__14258\,
            I => \N__14055\
        );

    \I__3312\ : ClkMux
    port map (
            O => \N__14257\,
            I => \N__14055\
        );

    \I__3311\ : ClkMux
    port map (
            O => \N__14256\,
            I => \N__14055\
        );

    \I__3310\ : ClkMux
    port map (
            O => \N__14255\,
            I => \N__14055\
        );

    \I__3309\ : ClkMux
    port map (
            O => \N__14254\,
            I => \N__14055\
        );

    \I__3308\ : ClkMux
    port map (
            O => \N__14253\,
            I => \N__14055\
        );

    \I__3307\ : ClkMux
    port map (
            O => \N__14252\,
            I => \N__14055\
        );

    \I__3306\ : ClkMux
    port map (
            O => \N__14251\,
            I => \N__14055\
        );

    \I__3305\ : ClkMux
    port map (
            O => \N__14250\,
            I => \N__14055\
        );

    \I__3304\ : ClkMux
    port map (
            O => \N__14249\,
            I => \N__14055\
        );

    \I__3303\ : ClkMux
    port map (
            O => \N__14248\,
            I => \N__14055\
        );

    \I__3302\ : ClkMux
    port map (
            O => \N__14247\,
            I => \N__14055\
        );

    \I__3301\ : ClkMux
    port map (
            O => \N__14246\,
            I => \N__14055\
        );

    \I__3300\ : ClkMux
    port map (
            O => \N__14245\,
            I => \N__14055\
        );

    \I__3299\ : ClkMux
    port map (
            O => \N__14244\,
            I => \N__14055\
        );

    \I__3298\ : ClkMux
    port map (
            O => \N__14243\,
            I => \N__14055\
        );

    \I__3297\ : ClkMux
    port map (
            O => \N__14242\,
            I => \N__14055\
        );

    \I__3296\ : ClkMux
    port map (
            O => \N__14241\,
            I => \N__14055\
        );

    \I__3295\ : ClkMux
    port map (
            O => \N__14240\,
            I => \N__14055\
        );

    \I__3294\ : ClkMux
    port map (
            O => \N__14239\,
            I => \N__14055\
        );

    \I__3293\ : ClkMux
    port map (
            O => \N__14238\,
            I => \N__14055\
        );

    \I__3292\ : ClkMux
    port map (
            O => \N__14237\,
            I => \N__14055\
        );

    \I__3291\ : ClkMux
    port map (
            O => \N__14236\,
            I => \N__14055\
        );

    \I__3290\ : ClkMux
    port map (
            O => \N__14235\,
            I => \N__14055\
        );

    \I__3289\ : ClkMux
    port map (
            O => \N__14234\,
            I => \N__14055\
        );

    \I__3288\ : ClkMux
    port map (
            O => \N__14233\,
            I => \N__14055\
        );

    \I__3287\ : ClkMux
    port map (
            O => \N__14232\,
            I => \N__14055\
        );

    \I__3286\ : ClkMux
    port map (
            O => \N__14231\,
            I => \N__14055\
        );

    \I__3285\ : ClkMux
    port map (
            O => \N__14230\,
            I => \N__14055\
        );

    \I__3284\ : ClkMux
    port map (
            O => \N__14229\,
            I => \N__14055\
        );

    \I__3283\ : ClkMux
    port map (
            O => \N__14228\,
            I => \N__14055\
        );

    \I__3282\ : ClkMux
    port map (
            O => \N__14227\,
            I => \N__14055\
        );

    \I__3281\ : ClkMux
    port map (
            O => \N__14226\,
            I => \N__14055\
        );

    \I__3280\ : ClkMux
    port map (
            O => \N__14225\,
            I => \N__14055\
        );

    \I__3279\ : ClkMux
    port map (
            O => \N__14224\,
            I => \N__14055\
        );

    \I__3278\ : ClkMux
    port map (
            O => \N__14223\,
            I => \N__14055\
        );

    \I__3277\ : ClkMux
    port map (
            O => \N__14222\,
            I => \N__14055\
        );

    \I__3276\ : ClkMux
    port map (
            O => \N__14221\,
            I => \N__14055\
        );

    \I__3275\ : ClkMux
    port map (
            O => \N__14220\,
            I => \N__14055\
        );

    \I__3274\ : ClkMux
    port map (
            O => \N__14219\,
            I => \N__14055\
        );

    \I__3273\ : ClkMux
    port map (
            O => \N__14218\,
            I => \N__14055\
        );

    \I__3272\ : ClkMux
    port map (
            O => \N__14217\,
            I => \N__14055\
        );

    \I__3271\ : ClkMux
    port map (
            O => \N__14216\,
            I => \N__14055\
        );

    \I__3270\ : ClkMux
    port map (
            O => \N__14215\,
            I => \N__14055\
        );

    \I__3269\ : ClkMux
    port map (
            O => \N__14214\,
            I => \N__14055\
        );

    \I__3268\ : ClkMux
    port map (
            O => \N__14213\,
            I => \N__14055\
        );

    \I__3267\ : ClkMux
    port map (
            O => \N__14212\,
            I => \N__14055\
        );

    \I__3266\ : ClkMux
    port map (
            O => \N__14211\,
            I => \N__14055\
        );

    \I__3265\ : ClkMux
    port map (
            O => \N__14210\,
            I => \N__14055\
        );

    \I__3264\ : ClkMux
    port map (
            O => \N__14209\,
            I => \N__14055\
        );

    \I__3263\ : ClkMux
    port map (
            O => \N__14208\,
            I => \N__14055\
        );

    \I__3262\ : ClkMux
    port map (
            O => \N__14207\,
            I => \N__14055\
        );

    \I__3261\ : ClkMux
    port map (
            O => \N__14206\,
            I => \N__14055\
        );

    \I__3260\ : ClkMux
    port map (
            O => \N__14205\,
            I => \N__14055\
        );

    \I__3259\ : ClkMux
    port map (
            O => \N__14204\,
            I => \N__14055\
        );

    \I__3258\ : GlobalMux
    port map (
            O => \N__14055\,
            I => \N__14052\
        );

    \I__3257\ : gio2CtrlBuf
    port map (
            O => \N__14052\,
            I => \CLK_c_g\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14046\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__14046\,
            I => \display2.prescaler_2_15\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__14043\,
            I => \N__14039\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \N__14033\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14023\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14023\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14023\
        );

    \I__3249\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14020\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14015\
        );

    \I__3247\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14015\
        );

    \I__3246\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14010\
        );

    \I__3245\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14010\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14023\,
            I => \N__14007\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__14020\,
            I => \display2.prescaler8_21\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__14015\,
            I => \display2.prescaler8_21\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__14010\,
            I => \display2.prescaler8_21\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__14007\,
            I => \display2.prescaler8_21\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__13998\,
            I => \display2.prescaler8_17_cascade_\
        );

    \I__3238\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13985\
        );

    \I__3237\ : InMux
    port map (
            O => \N__13994\,
            I => \N__13985\
        );

    \I__3236\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13973\
        );

    \I__3235\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13973\
        );

    \I__3234\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13973\
        );

    \I__3233\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13973\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__13985\,
            I => \N__13970\
        );

    \I__3231\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13963\
        );

    \I__3230\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13963\
        );

    \I__3229\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13963\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__13973\,
            I => \N__13960\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__13970\,
            I => \display2.prescaler8_16\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__13963\,
            I => \display2.prescaler8_16\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__13960\,
            I => \display2.prescaler8_16\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__13953\,
            I => \N__13949\
        );

    \I__3223\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13946\
        );

    \I__3222\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13943\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__13946\,
            I => \display2.prescalerZ0Z_15\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__13943\,
            I => \display2.prescalerZ0Z_15\
        );

    \I__3219\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__13935\,
            I => \N__13932\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__13932\,
            I => \N__13929\
        );

    \I__3216\ : Sp12to4
    port map (
            O => \N__13929\,
            I => \N__13926\
        );

    \I__3215\ : Span12Mux_h
    port map (
            O => \N__13926\,
            I => \N__13923\
        );

    \I__3214\ : Span12Mux_v
    port map (
            O => \N__13923\,
            I => \N__13920\
        );

    \I__3213\ : Odrv12
    port map (
            O => \N__13920\,
            I => switch_up_c
        );

    \I__3212\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13914\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__13914\,
            I => \N__13911\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__13911\,
            I => \N__13908\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__13908\,
            I => \N__13905\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__13905\,
            I => \N__13902\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__13902\,
            I => \d1.syncZ0Z_0\
        );

    \I__3206\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13893\
        );

    \I__3205\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13889\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__13897\,
            I => \N__13886\
        );

    \I__3203\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13882\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__13893\,
            I => \N__13879\
        );

    \I__3201\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13876\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__13889\,
            I => \N__13873\
        );

    \I__3199\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13868\
        );

    \I__3198\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13868\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__13882\,
            I => \N__13863\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__13879\,
            I => \N__13859\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__13876\,
            I => \N__13856\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__13873\,
            I => \N__13851\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__13868\,
            I => \N__13851\
        );

    \I__3192\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13845\
        );

    \I__3191\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13842\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__13863\,
            I => \N__13838\
        );

    \I__3189\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13835\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__13859\,
            I => \N__13828\
        );

    \I__3187\ : Span4Mux_v
    port map (
            O => \N__13856\,
            I => \N__13828\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__13851\,
            I => \N__13828\
        );

    \I__3185\ : InMux
    port map (
            O => \N__13850\,
            I => \N__13825\
        );

    \I__3184\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13820\
        );

    \I__3183\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13820\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__13845\,
            I => \N__13817\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__13842\,
            I => \N__13814\
        );

    \I__3180\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13811\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__13838\,
            I => \minsZ0Z_3\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__13835\,
            I => \minsZ0Z_3\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__13828\,
            I => \minsZ0Z_3\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__13825\,
            I => \minsZ0Z_3\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__13820\,
            I => \minsZ0Z_3\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__13817\,
            I => \minsZ0Z_3\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__13814\,
            I => \minsZ0Z_3\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__13811\,
            I => \minsZ0Z_3\
        );

    \I__3171\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13791\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__13791\,
            I => \N__13785\
        );

    \I__3169\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13782\
        );

    \I__3168\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13777\
        );

    \I__3167\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13773\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__13785\,
            I => \N__13769\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__13782\,
            I => \N__13766\
        );

    \I__3164\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13761\
        );

    \I__3163\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13758\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__13777\,
            I => \N__13752\
        );

    \I__3161\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13749\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__13773\,
            I => \N__13744\
        );

    \I__3159\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13741\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__13769\,
            I => \N__13736\
        );

    \I__3157\ : Span4Mux_v
    port map (
            O => \N__13766\,
            I => \N__13736\
        );

    \I__3156\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13731\
        );

    \I__3155\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13731\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13728\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__13758\,
            I => \N__13725\
        );

    \I__3152\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13720\
        );

    \I__3151\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13720\
        );

    \I__3150\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13717\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__13752\,
            I => \N__13714\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__13749\,
            I => \N__13711\
        );

    \I__3147\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13706\
        );

    \I__3146\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13706\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__13744\,
            I => \minsZ0Z_2\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__13741\,
            I => \minsZ0Z_2\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__13736\,
            I => \minsZ0Z_2\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__13731\,
            I => \minsZ0Z_2\
        );

    \I__3141\ : Odrv12
    port map (
            O => \N__13728\,
            I => \minsZ0Z_2\
        );

    \I__3140\ : Odrv12
    port map (
            O => \N__13725\,
            I => \minsZ0Z_2\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__13720\,
            I => \minsZ0Z_2\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__13717\,
            I => \minsZ0Z_2\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__13714\,
            I => \minsZ0Z_2\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__13711\,
            I => \minsZ0Z_2\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__13706\,
            I => \minsZ0Z_2\
        );

    \I__3134\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13676\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__13682\,
            I => \N__13672\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \N__13667\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__13680\,
            I => \N__13664\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__13679\,
            I => \N__13661\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__13676\,
            I => \N__13658\
        );

    \I__3128\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13655\
        );

    \I__3127\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13652\
        );

    \I__3126\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13647\
        );

    \I__3125\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13641\
        );

    \I__3124\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13641\
        );

    \I__3123\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13638\
        );

    \I__3122\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13635\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__13658\,
            I => \N__13626\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__13655\,
            I => \N__13626\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13623\
        );

    \I__3118\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13618\
        );

    \I__3117\ : InMux
    port map (
            O => \N__13650\,
            I => \N__13618\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__13647\,
            I => \N__13615\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__13646\,
            I => \N__13611\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__13641\,
            I => \N__13604\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__13638\,
            I => \N__13604\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13604\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__13634\,
            I => \N__13601\
        );

    \I__3110\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13598\
        );

    \I__3109\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13595\
        );

    \I__3108\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13592\
        );

    \I__3107\ : Span4Mux_h
    port map (
            O => \N__13626\,
            I => \N__13585\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__13623\,
            I => \N__13585\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__13618\,
            I => \N__13585\
        );

    \I__3104\ : Span4Mux_h
    port map (
            O => \N__13615\,
            I => \N__13582\
        );

    \I__3103\ : InMux
    port map (
            O => \N__13614\,
            I => \N__13577\
        );

    \I__3102\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13577\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__13604\,
            I => \N__13574\
        );

    \I__3100\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13571\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__13598\,
            I => \minsZ0Z_1\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__13595\,
            I => \minsZ0Z_1\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__13592\,
            I => \minsZ0Z_1\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__13585\,
            I => \minsZ0Z_1\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__13582\,
            I => \minsZ0Z_1\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__13577\,
            I => \minsZ0Z_1\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__13574\,
            I => \minsZ0Z_1\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__13571\,
            I => \minsZ0Z_1\
        );

    \I__3091\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13551\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__13551\,
            I => \N__13539\
        );

    \I__3089\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13536\
        );

    \I__3088\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13532\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__13548\,
            I => \N__13529\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__13547\,
            I => \N__13526\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__13546\,
            I => \N__13523\
        );

    \I__3084\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13518\
        );

    \I__3083\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13518\
        );

    \I__3082\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13515\
        );

    \I__3081\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13512\
        );

    \I__3080\ : Span4Mux_v
    port map (
            O => \N__13539\,
            I => \N__13507\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__13536\,
            I => \N__13504\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__13535\,
            I => \N__13500\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13496\
        );

    \I__3076\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13493\
        );

    \I__3075\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13490\
        );

    \I__3074\ : InMux
    port map (
            O => \N__13523\,
            I => \N__13484\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__13518\,
            I => \N__13481\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13476\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13512\,
            I => \N__13476\
        );

    \I__3070\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13473\
        );

    \I__3069\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13470\
        );

    \I__3068\ : Span4Mux_h
    port map (
            O => \N__13507\,
            I => \N__13465\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__13504\,
            I => \N__13465\
        );

    \I__3066\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13458\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13458\
        );

    \I__3064\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13458\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__13496\,
            I => \N__13453\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__13493\,
            I => \N__13453\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__13490\,
            I => \N__13450\
        );

    \I__3060\ : InMux
    port map (
            O => \N__13489\,
            I => \N__13445\
        );

    \I__3059\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13445\
        );

    \I__3058\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13442\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13435\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__13481\,
            I => \N__13435\
        );

    \I__3055\ : Span4Mux_h
    port map (
            O => \N__13476\,
            I => \N__13435\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__13473\,
            I => \minsZ0Z_0\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__13470\,
            I => \minsZ0Z_0\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__13465\,
            I => \minsZ0Z_0\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__13458\,
            I => \minsZ0Z_0\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__13453\,
            I => \minsZ0Z_0\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__13450\,
            I => \minsZ0Z_0\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__13445\,
            I => \minsZ0Z_0\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__13442\,
            I => \minsZ0Z_0\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__13435\,
            I => \minsZ0Z_0\
        );

    \I__3045\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13413\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__13413\,
            I => \N__13407\
        );

    \I__3043\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13402\
        );

    \I__3042\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13402\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__13410\,
            I => \N__13397\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__13407\,
            I => \N__13394\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__13402\,
            I => \N__13391\
        );

    \I__3038\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13386\
        );

    \I__3037\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13386\
        );

    \I__3036\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13383\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__13394\,
            I => \display2.digit_posnZ0\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__13391\,
            I => \display2.digit_posnZ0\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__13386\,
            I => \display2.digit_posnZ0\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__13383\,
            I => \display2.digit_posnZ0\
        );

    \I__3031\ : IoInMux
    port map (
            O => \N__13374\,
            I => \N__13371\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__13371\,
            I => \N__13368\
        );

    \I__3029\ : IoSpan4Mux
    port map (
            O => \N__13368\,
            I => \N__13365\
        );

    \I__3028\ : Span4Mux_s2_h
    port map (
            O => \N__13365\,
            I => \N__13362\
        );

    \I__3027\ : Sp12to4
    port map (
            O => \N__13362\,
            I => \N__13359\
        );

    \I__3026\ : Span12Mux_s11_h
    port map (
            O => \N__13359\,
            I => \N__13356\
        );

    \I__3025\ : Odrv12
    port map (
            O => \N__13356\,
            I => \DIGIT_c_1\
        );

    \I__3024\ : CEMux
    port map (
            O => \N__13353\,
            I => \N__13350\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__13350\,
            I => \N__13347\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__13347\,
            I => \N__13340\
        );

    \I__3021\ : InMux
    port map (
            O => \N__13346\,
            I => \N__13335\
        );

    \I__3020\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13335\
        );

    \I__3019\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13330\
        );

    \I__3018\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13330\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__13340\,
            I => \display2.prescaler8\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13335\,
            I => \display2.prescaler8\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__13330\,
            I => \display2.prescaler8\
        );

    \I__3014\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13320\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__3012\ : Span12Mux_h
    port map (
            O => \N__13317\,
            I => \N__13314\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__13314\,
            I => switch_start_stop_c
        );

    \I__3010\ : InMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__3008\ : Span12Mux_v
    port map (
            O => \N__13305\,
            I => \N__13302\
        );

    \I__3007\ : Odrv12
    port map (
            O => \N__13302\,
            I => \d4.syncZ0Z_0\
        );

    \I__3006\ : IoInMux
    port map (
            O => \N__13299\,
            I => \N__13296\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__13296\,
            I => \N__13293\
        );

    \I__3004\ : Span4Mux_s2_h
    port map (
            O => \N__13293\,
            I => \N__13290\
        );

    \I__3003\ : Span4Mux_v
    port map (
            O => \N__13290\,
            I => \N__13287\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__13287\,
            I => \SEG2_c_0\
        );

    \I__3001\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13280\
        );

    \I__3000\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13277\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__13280\,
            I => \N__13274\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__13277\,
            I => \display2.prescalerZ0Z_12\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__13274\,
            I => \display2.prescalerZ0Z_12\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13265\
        );

    \I__2995\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13262\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__13265\,
            I => \display2.prescalerZ0Z_10\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__13262\,
            I => \display2.prescalerZ0Z_10\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__13257\,
            I => \N__13254\
        );

    \I__2991\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13250\
        );

    \I__2990\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13247\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13244\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__13247\,
            I => \display2.prescalerZ0Z_13\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__13244\,
            I => \display2.prescalerZ0Z_13\
        );

    \I__2986\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13235\
        );

    \I__2985\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13232\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__13235\,
            I => \display2.prescalerZ0Z_11\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13232\,
            I => \display2.prescalerZ0Z_11\
        );

    \I__2982\ : InMux
    port map (
            O => \N__13227\,
            I => \N__13224\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__13221\,
            I => \display2.prescaler8_15\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__13218\,
            I => \display2.prescaler8_12_cascade_\
        );

    \I__2978\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13212\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__13212\,
            I => \display2.prescaler8_13\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__13209\,
            I => \display2.prescaler8_21_cascade_\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__13206\,
            I => \N__13201\
        );

    \I__2974\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13198\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13195\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13192\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__13198\,
            I => \display2.prescalerZ0Z_1\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__13195\,
            I => \display2.prescalerZ0Z_1\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__13192\,
            I => \display2.prescalerZ0Z_1\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__13182\,
            I => \display2.prescaler8_14\
        );

    \I__2966\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__13176\,
            I => \display2.prescaler_2_9\
        );

    \I__2964\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13169\
        );

    \I__2963\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13166\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__13169\,
            I => \display2.prescalerZ0Z_9\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__13166\,
            I => \display2.prescalerZ0Z_9\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13158\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__13158\,
            I => \display2.prescaler_2_14\
        );

    \I__2958\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13151\
        );

    \I__2957\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13148\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__13151\,
            I => \display2.prescalerZ0Z_14\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__13148\,
            I => \display2.prescalerZ0Z_14\
        );

    \I__2954\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13139\
        );

    \I__2953\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__13139\,
            I => \display2.prescalerZ0Z_17\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__13136\,
            I => \display2.prescalerZ0Z_17\
        );

    \I__2950\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13127\
        );

    \I__2949\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13124\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__13127\,
            I => \display2.prescalerZ0Z_16\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__13124\,
            I => \display2.prescalerZ0Z_16\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \N__13115\
        );

    \I__2945\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13112\
        );

    \I__2944\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13109\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__13112\,
            I => \display2.prescalerZ0Z_18\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__13109\,
            I => \display2.prescalerZ0Z_18\
        );

    \I__2941\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13096\
        );

    \I__2940\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13096\
        );

    \I__2939\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13093\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13090\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__13096\,
            I => \display2.prescalerZ0Z_0\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__13093\,
            I => \display2.prescalerZ0Z_0\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__13090\,
            I => \display2.prescalerZ0Z_0\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__13083\,
            I => \N__13078\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__13082\,
            I => \N__13075\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__13081\,
            I => \N__13070\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13061\
        );

    \I__2930\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13061\
        );

    \I__2929\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13061\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \N__13058\
        );

    \I__2927\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13054\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13049\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13049\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13046\
        );

    \I__2923\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13041\
        );

    \I__2922\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13041\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__13054\,
            I => \display2.prescaler8_17\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__13049\,
            I => \display2.prescaler8_17\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__13046\,
            I => \display2.prescaler8_17\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__13041\,
            I => \display2.prescaler8_17\
        );

    \I__2917\ : InMux
    port map (
            O => \N__13032\,
            I => \display2.prescaler_2_cry_18\
        );

    \I__2916\ : InMux
    port map (
            O => \N__13029\,
            I => \display2.prescaler_2_cry_19\
        );

    \I__2915\ : InMux
    port map (
            O => \N__13026\,
            I => \display2.prescaler_2_cry_20\
        );

    \I__2914\ : InMux
    port map (
            O => \N__13023\,
            I => \display2.prescaler_2_cry_21\
        );

    \I__2913\ : InMux
    port map (
            O => \N__13020\,
            I => \display2.prescaler_2_cry_22\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__13017\,
            I => \N__13013\
        );

    \I__2911\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13010\
        );

    \I__2910\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13007\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__13010\,
            I => \display2.prescalerZ0Z_23\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__13007\,
            I => \display2.prescalerZ0Z_23\
        );

    \I__2907\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12996\
        );

    \I__2906\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12996\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__12996\,
            I => \display2.prescalerZ0Z_21\
        );

    \I__2904\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12987\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12987\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__12987\,
            I => \display2.prescalerZ0Z_20\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__12984\,
            I => \N__12980\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \N__12977\
        );

    \I__2899\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12972\
        );

    \I__2898\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12972\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__12972\,
            I => \display2.prescalerZ0Z_22\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__12969\,
            I => \N__12966\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12960\
        );

    \I__2894\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12960\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__12960\,
            I => \display2.prescalerZ0Z_19\
        );

    \I__2892\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12953\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12950\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__12953\,
            I => \display2.prescalerZ0Z_5\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__12950\,
            I => \display2.prescalerZ0Z_5\
        );

    \I__2888\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12941\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12938\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__12941\,
            I => \display2.prescalerZ0Z_3\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__12938\,
            I => \display2.prescalerZ0Z_3\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__12933\,
            I => \N__12929\
        );

    \I__2883\ : InMux
    port map (
            O => \N__12932\,
            I => \N__12926\
        );

    \I__2882\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12923\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__12926\,
            I => \display2.prescalerZ0Z_7\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__12923\,
            I => \display2.prescalerZ0Z_7\
        );

    \I__2879\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12914\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12911\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__12914\,
            I => \display2.prescalerZ0Z_2\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__12911\,
            I => \display2.prescalerZ0Z_2\
        );

    \I__2875\ : InMux
    port map (
            O => \N__12906\,
            I => \display2.prescaler_2_cry_9\
        );

    \I__2874\ : InMux
    port map (
            O => \N__12903\,
            I => \display2.prescaler_2_cry_10\
        );

    \I__2873\ : InMux
    port map (
            O => \N__12900\,
            I => \display2.prescaler_2_cry_11\
        );

    \I__2872\ : InMux
    port map (
            O => \N__12897\,
            I => \display2.prescaler_2_cry_12\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12894\,
            I => \display2.prescaler_2_cry_13\
        );

    \I__2870\ : InMux
    port map (
            O => \N__12891\,
            I => \display2.prescaler_2_cry_14\
        );

    \I__2869\ : InMux
    port map (
            O => \N__12888\,
            I => \display2.prescaler_2_cry_15\
        );

    \I__2868\ : InMux
    port map (
            O => \N__12885\,
            I => \bfn_14_14_0_\
        );

    \I__2867\ : InMux
    port map (
            O => \N__12882\,
            I => \display2.prescaler_2_cry_17\
        );

    \I__2866\ : InMux
    port map (
            O => \N__12879\,
            I => \display2.prescaler_2_cry_1\
        );

    \I__2865\ : InMux
    port map (
            O => \N__12876\,
            I => \display2.prescaler_2_cry_2\
        );

    \I__2864\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12869\
        );

    \I__2863\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12866\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__12869\,
            I => \display2.prescalerZ0Z_4\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__12866\,
            I => \display2.prescalerZ0Z_4\
        );

    \I__2860\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12858\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__12858\,
            I => \display2.prescaler_2_4\
        );

    \I__2858\ : InMux
    port map (
            O => \N__12855\,
            I => \display2.prescaler_2_cry_3\
        );

    \I__2857\ : InMux
    port map (
            O => \N__12852\,
            I => \display2.prescaler_2_cry_4\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12845\
        );

    \I__2855\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12842\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__12845\,
            I => \display2.prescalerZ0Z_6\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12842\,
            I => \display2.prescalerZ0Z_6\
        );

    \I__2852\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12834\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__12834\,
            I => \display2.prescaler_2_6\
        );

    \I__2850\ : InMux
    port map (
            O => \N__12831\,
            I => \display2.prescaler_2_cry_5\
        );

    \I__2849\ : InMux
    port map (
            O => \N__12828\,
            I => \display2.prescaler_2_cry_6\
        );

    \I__2848\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12821\
        );

    \I__2847\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12818\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__12821\,
            I => \display2.prescalerZ0Z_8\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__12818\,
            I => \display2.prescalerZ0Z_8\
        );

    \I__2844\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12810\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12810\,
            I => \display2.prescaler_2_8\
        );

    \I__2842\ : InMux
    port map (
            O => \N__12807\,
            I => \display2.prescaler_2_cry_7\
        );

    \I__2841\ : InMux
    port map (
            O => \N__12804\,
            I => \bfn_14_13_0_\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__12801\,
            I => \N__12792\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__12800\,
            I => \N__12786\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__12799\,
            I => \N__12781\
        );

    \I__2837\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12778\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__12797\,
            I => \N__12775\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__12796\,
            I => \N__12771\
        );

    \I__2834\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12763\
        );

    \I__2833\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12763\
        );

    \I__2832\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12763\
        );

    \I__2831\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12760\
        );

    \I__2830\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12756\
        );

    \I__2829\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12753\
        );

    \I__2828\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12750\
        );

    \I__2827\ : InMux
    port map (
            O => \N__12784\,
            I => \N__12745\
        );

    \I__2826\ : InMux
    port map (
            O => \N__12781\,
            I => \N__12742\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__12778\,
            I => \N__12739\
        );

    \I__2824\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12736\
        );

    \I__2823\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12733\
        );

    \I__2822\ : InMux
    port map (
            O => \N__12771\,
            I => \N__12726\
        );

    \I__2821\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12726\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12723\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__12760\,
            I => \N__12720\
        );

    \I__2818\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12717\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__12756\,
            I => \N__12709\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__12753\,
            I => \N__12709\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__12750\,
            I => \N__12709\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12706\
        );

    \I__2813\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12703\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__12745\,
            I => \N__12700\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__12742\,
            I => \N__12695\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__12739\,
            I => \N__12695\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__12736\,
            I => \N__12690\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__12733\,
            I => \N__12690\
        );

    \I__2807\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12685\
        );

    \I__2806\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12685\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__12726\,
            I => \N__12681\
        );

    \I__2804\ : Span4Mux_h
    port map (
            O => \N__12723\,
            I => \N__12676\
        );

    \I__2803\ : Span4Mux_h
    port map (
            O => \N__12720\,
            I => \N__12676\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12717\,
            I => \N__12673\
        );

    \I__2801\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12670\
        );

    \I__2800\ : Span4Mux_v
    port map (
            O => \N__12709\,
            I => \N__12667\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__12706\,
            I => \N__12656\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12703\,
            I => \N__12656\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__12700\,
            I => \N__12656\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__12695\,
            I => \N__12656\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__12690\,
            I => \N__12656\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__12685\,
            I => \N__12653\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12684\,
            I => \N__12650\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__12681\,
            I => \N__12647\
        );

    \I__2791\ : Span4Mux_v
    port map (
            O => \N__12676\,
            I => \N__12642\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__12673\,
            I => \N__12642\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__12670\,
            I => \stateZ0Z_0\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__12667\,
            I => \stateZ0Z_0\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__12656\,
            I => \stateZ0Z_0\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__12653\,
            I => \stateZ0Z_0\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__12650\,
            I => \stateZ0Z_0\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__12647\,
            I => \stateZ0Z_0\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__12642\,
            I => \stateZ0Z_0\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__12627\,
            I => \d2_g0_1_cascade_\
        );

    \I__2781\ : InMux
    port map (
            O => \N__12624\,
            I => \N__12621\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__12621\,
            I => \d1.g2_i_a5_1Z0Z_3\
        );

    \I__2779\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12614\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12611\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__12614\,
            I => \N__12606\
        );

    \I__2776\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12603\
        );

    \I__2775\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12600\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12597\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__12606\,
            I => \N__12592\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__12603\,
            I => \N__12592\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__12600\,
            I => \N__12587\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__12597\,
            I => \N__12587\
        );

    \I__2769\ : Span4Mux_h
    port map (
            O => \N__12592\,
            I => \N__12584\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__12587\,
            I => \N__12581\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__12584\,
            I => \d3.syncZ0Z_1\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__12581\,
            I => \d3.syncZ0Z_1\
        );

    \I__2765\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12572\
        );

    \I__2764\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12569\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12564\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__12569\,
            I => \N__12561\
        );

    \I__2761\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12558\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12555\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__12564\,
            I => \N__12552\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__12561\,
            I => \d3.stateZ0\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__12558\,
            I => \d3.stateZ0\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12555\,
            I => \d3.stateZ0\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__12552\,
            I => \d3.stateZ0\
        );

    \I__2754\ : IoInMux
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12537\
        );

    \I__2752\ : Span4Mux_s2_h
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__2750\ : Span4Mux_h
    port map (
            O => \N__12531\,
            I => \N__12528\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__12528\,
            I => \N__12525\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__12525\,
            I => \d3.idle_i\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__2746\ : InMux
    port map (
            O => \N__12519\,
            I => \N__12516\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__12516\,
            I => \N__12513\
        );

    \I__2744\ : Span4Mux_v
    port map (
            O => \N__12513\,
            I => \N__12510\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__12510\,
            I => \d1.g0_1_0Z0Z_0\
        );

    \I__2742\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12502\
        );

    \I__2741\ : InMux
    port map (
            O => \N__12506\,
            I => \N__12499\
        );

    \I__2740\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12496\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12502\,
            I => \N__12491\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12499\,
            I => \N__12485\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12485\
        );

    \I__2736\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12482\
        );

    \I__2735\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12479\
        );

    \I__2734\ : Span12Mux_h
    port map (
            O => \N__12491\,
            I => \N__12476\
        );

    \I__2733\ : InMux
    port map (
            O => \N__12490\,
            I => \N__12473\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__12485\,
            I => \N__12468\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__12482\,
            I => \N__12468\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__12479\,
            I => \N__12465\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__12476\,
            I => \ten_secsZ0Z_1\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__12473\,
            I => \ten_secsZ0Z_1\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__12468\,
            I => \ten_secsZ0Z_1\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__12465\,
            I => \ten_secsZ0Z_1\
        );

    \I__2725\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12453\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__12453\,
            I => \N__12446\
        );

    \I__2723\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12443\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12440\
        );

    \I__2721\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12437\
        );

    \I__2720\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12433\
        );

    \I__2719\ : Span4Mux_h
    port map (
            O => \N__12446\,
            I => \N__12430\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__12443\,
            I => \N__12426\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__12440\,
            I => \N__12421\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12421\
        );

    \I__2715\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12418\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__12433\,
            I => \N__12415\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__12430\,
            I => \N__12412\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12429\,
            I => \N__12409\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__12426\,
            I => \N__12404\
        );

    \I__2710\ : Span4Mux_v
    port map (
            O => \N__12421\,
            I => \N__12404\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__12418\,
            I => \N__12399\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__12415\,
            I => \N__12399\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__12412\,
            I => \ten_secsZ0Z_0\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__12409\,
            I => \ten_secsZ0Z_0\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__12404\,
            I => \ten_secsZ0Z_0\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__12399\,
            I => \ten_secsZ0Z_0\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__12390\,
            I => \N__12387\
        );

    \I__2702\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12384\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__12381\,
            I => \N__12378\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__12375\,
            I => \BNC1\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12367\
        );

    \I__2696\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12362\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12362\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__12367\,
            I => \d2.countZ0Z_9\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__12362\,
            I => \d2.countZ0Z_9\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__12357\,
            I => \N__12353\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12349\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12345\
        );

    \I__2689\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12342\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__12349\,
            I => \N__12338\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__12348\,
            I => \N__12334\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12345\,
            I => \N__12331\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12328\
        );

    \I__2684\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12323\
        );

    \I__2683\ : Span4Mux_h
    port map (
            O => \N__12338\,
            I => \N__12320\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12315\
        );

    \I__2681\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12315\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__12331\,
            I => \N__12310\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__12328\,
            I => \N__12310\
        );

    \I__2678\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12305\
        );

    \I__2677\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12305\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__12323\,
            I => d2_count_16
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__12320\,
            I => d2_count_16
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12315\,
            I => d2_count_16
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__12310\,
            I => d2_count_16
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__12305\,
            I => d2_count_16
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__12294\,
            I => \N__12289\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__12293\,
            I => \N__12286\
        );

    \I__2669\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12283\
        );

    \I__2668\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12278\
        );

    \I__2667\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12278\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__12283\,
            I => \d2.countZ0Z_10\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__12278\,
            I => \d2.countZ0Z_10\
        );

    \I__2664\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12268\
        );

    \I__2663\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__2662\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12263\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__12268\,
            I => \d2.countZ0Z_7\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__12263\,
            I => \d2.countZ0Z_7\
        );

    \I__2659\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12255\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__12255\,
            I => \N__12252\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__12252\,
            I => \d2.g0_0_13\
        );

    \I__2656\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12239\
        );

    \I__2655\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12236\
        );

    \I__2654\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12233\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12228\
        );

    \I__2652\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12228\
        );

    \I__2651\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12223\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12223\
        );

    \I__2649\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12220\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__12239\,
            I => \N__12217\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__12236\,
            I => d2_count_3
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__12233\,
            I => d2_count_3
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__12228\,
            I => d2_count_3
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__12223\,
            I => d2_count_3
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__12220\,
            I => d2_count_3
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__12217\,
            I => d2_count_3
        );

    \I__2641\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12201\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__12201\,
            I => \d1.g2_8_2\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__12198\,
            I => \N__12194\
        );

    \I__2638\ : InMux
    port map (
            O => \N__12197\,
            I => \N__12190\
        );

    \I__2637\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12187\
        );

    \I__2636\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12184\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__12190\,
            I => \d2.countZ0Z_12\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__12187\,
            I => \d2.countZ0Z_12\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__12184\,
            I => \d2.countZ0Z_12\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__12177\,
            I => \N__12172\
        );

    \I__2631\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12169\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12166\
        );

    \I__2629\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12163\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__12169\,
            I => \d2.countZ0Z_13\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__12166\,
            I => \d2.countZ0Z_13\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__12163\,
            I => \d2.countZ0Z_13\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \N__12152\
        );

    \I__2624\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12148\
        );

    \I__2623\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12145\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12142\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__12148\,
            I => \d2.countZ0Z_14\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__12145\,
            I => \d2.countZ0Z_14\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__12142\,
            I => \d2.countZ0Z_14\
        );

    \I__2618\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12131\
        );

    \I__2617\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12127\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12124\
        );

    \I__2615\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12121\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__12127\,
            I => \d2.countZ0Z_11\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__12124\,
            I => \d2.countZ0Z_11\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__12121\,
            I => \d2.countZ0Z_11\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12110\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12106\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__12110\,
            I => \N__12103\
        );

    \I__2608\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12097\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12106\,
            I => \N__12093\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__12103\,
            I => \N__12090\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__12102\,
            I => \N__12087\
        );

    \I__2604\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12082\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12100\,
            I => \N__12082\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__12097\,
            I => \N__12079\
        );

    \I__2601\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12076\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__12093\,
            I => \N__12071\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__12090\,
            I => \N__12071\
        );

    \I__2598\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12068\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12063\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__12079\,
            I => \N__12063\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__12076\,
            I => d2_trans_up_1_15_7
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__12071\,
            I => d2_trans_up_1_15_7
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__12068\,
            I => d2_trans_up_1_15_7
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__12063\,
            I => d2_trans_up_1_15_7
        );

    \I__2591\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12051\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__12051\,
            I => \d1.g2_i_a5_1Z0Z_6\
        );

    \I__2589\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12039\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__12046\,
            I => \N__12036\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__12045\,
            I => \N__12033\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__12042\,
            I => \N__12029\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12026\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12022\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12019\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__12032\,
            I => \N__12014\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__12029\,
            I => \N__12009\
        );

    \I__2579\ : Span4Mux_h
    port map (
            O => \N__12026\,
            I => \N__12009\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12025\,
            I => \N__12006\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__12001\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__12001\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12018\,
            I => \N__11994\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12017\,
            I => \N__11994\
        );

    \I__2573\ : InMux
    port map (
            O => \N__12014\,
            I => \N__11994\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__12009\,
            I => d2_sync_1
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__12006\,
            I => d2_sync_1
        );

    \I__2570\ : Odrv12
    port map (
            O => \N__12001\,
            I => d2_sync_1
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11994\,
            I => d2_sync_1
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__11985\,
            I => \N__11982\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11977\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11974\
        );

    \I__2565\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11969\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11964\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__11974\,
            I => \N__11964\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11959\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11959\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11969\,
            I => \N__11955\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__11964\,
            I => \N__11950\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11959\,
            I => \N__11950\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11946\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__11955\,
            I => \N__11940\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__11950\,
            I => \N__11940\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11933\
        );

    \I__2553\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11933\
        );

    \I__2552\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11933\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__11940\,
            I => d2_state
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__11933\,
            I => d2_state
        );

    \I__2549\ : IoInMux
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__11922\,
            I => \d2.idle_i\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11915\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__11915\,
            I => d2_g0_3
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__11912\,
            I => d2_g0_3
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__11907\,
            I => \d1.g0_1_0_a4Z0Z_4_cascade_\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11895\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11892\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11883\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11878\
        );

    \I__2537\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11873\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11873\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11870\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11895\,
            I => \N__11865\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11892\,
            I => \N__11865\
        );

    \I__2532\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11853\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11853\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11853\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11846\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11846\
        );

    \I__2527\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11846\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11843\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11838\
        );

    \I__2524\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11838\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11829\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11829\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__11870\,
            I => \N__11829\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__11865\,
            I => \N__11829\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11826\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11823\
        );

    \I__2517\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11818\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11818\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11815\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11810\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11846\,
            I => \N__11810\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__11843\,
            I => \N__11807\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11838\,
            I => \N__11804\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__11829\,
            I => \N__11801\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11826\,
            I => \N__11794\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__11823\,
            I => \N__11794\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__11818\,
            I => \N__11794\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__11815\,
            I => \N__11791\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__11810\,
            I => \N__11784\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__11807\,
            I => \N__11784\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__11804\,
            I => \N__11784\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__11801\,
            I => \stateZ0Z_1\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__11794\,
            I => \stateZ0Z_1\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__11791\,
            I => \stateZ0Z_1\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__11784\,
            I => \stateZ0Z_1\
        );

    \I__2498\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__2496\ : Odrv12
    port map (
            O => \N__11769\,
            I => \d1.g0_1_0_a4Z0Z_8\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__11766\,
            I => \N__11762\
        );

    \I__2494\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11754\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11754\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__11761\,
            I => \N__11748\
        );

    \I__2491\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11744\
        );

    \I__2490\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11741\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11738\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11735\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11728\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11728\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11728\
        );

    \I__2484\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11725\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11744\,
            I => d2_count_15
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11741\,
            I => d2_count_15
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__11738\,
            I => d2_count_15
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11735\,
            I => d2_count_15
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__11728\,
            I => d2_count_15
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__11725\,
            I => d2_count_15
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \N__11707\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__11711\,
            I => \N__11704\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11701\
        );

    \I__2474\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11698\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11691\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11701\,
            I => \N__11686\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11698\,
            I => \N__11686\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__11697\,
            I => \N__11681\
        );

    \I__2469\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11677\
        );

    \I__2468\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11674\
        );

    \I__2467\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11671\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__11691\,
            I => \N__11666\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__11686\,
            I => \N__11666\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11661\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11661\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11656\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11656\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__11677\,
            I => d2_count_2
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__11674\,
            I => d2_count_2
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__11671\,
            I => d2_count_2
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__11666\,
            I => d2_count_2
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11661\,
            I => d2_count_2
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__11656\,
            I => d2_count_2
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__11643\,
            I => \N__11640\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11635\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11629\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11629\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__11635\,
            I => \N__11623\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11617\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__11629\,
            I => \N__11614\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11609\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11609\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11605\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__11623\,
            I => \N__11602\
        );

    \I__2443\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11599\
        );

    \I__2442\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11594\
        );

    \I__2441\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11594\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__11617\,
            I => \N__11591\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__11614\,
            I => \N__11586\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11586\
        );

    \I__2437\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11583\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__11605\,
            I => d2_count_1
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__11602\,
            I => d2_count_1
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__11599\,
            I => d2_count_1
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__11594\,
            I => d2_count_1
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__11591\,
            I => d2_count_1
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__11586\,
            I => d2_count_1
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__11583\,
            I => d2_count_1
        );

    \I__2429\ : SRMux
    port map (
            O => \N__11568\,
            I => \N__11565\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11565\,
            I => \N__11561\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__11564\,
            I => \N__11558\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__11561\,
            I => \N__11555\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N__11552\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__11555\,
            I => \N__11548\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__11552\,
            I => \N__11545\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__11551\,
            I => \N__11542\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__11548\,
            I => \N__11538\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__11545\,
            I => \N__11535\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__11542\,
            I => \N__11532\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11529\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__11538\,
            I => mins_0_sqmuxa
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__11535\,
            I => mins_0_sqmuxa
        );

    \I__2415\ : Odrv12
    port map (
            O => \N__11532\,
            I => mins_0_sqmuxa
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__11529\,
            I => mins_0_sqmuxa
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11514\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__2410\ : Span4Mux_h
    port map (
            O => \N__11511\,
            I => \N__11508\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__11508\,
            I => \d1.g0_1_a5_0Z0Z_11\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11502\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__11499\,
            I => \N__11496\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__11496\,
            I => \d1.g2_12_1\
        );

    \I__2404\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11489\
        );

    \I__2403\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11485\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__11489\,
            I => \N__11481\
        );

    \I__2401\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11475\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__11485\,
            I => \N__11472\
        );

    \I__2399\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11469\
        );

    \I__2398\ : Span4Mux_h
    port map (
            O => \N__11481\,
            I => \N__11466\
        );

    \I__2397\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11459\
        );

    \I__2396\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11459\
        );

    \I__2395\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11459\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__11475\,
            I => d2_count_4
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__11472\,
            I => d2_count_4
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__11469\,
            I => d2_count_4
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__11466\,
            I => d2_count_4
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__11459\,
            I => d2_count_4
        );

    \I__2389\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11444\
        );

    \I__2388\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11441\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11435\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11431\
        );

    \I__2385\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11428\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11420\
        );

    \I__2383\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11420\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__11435\,
            I => \N__11417\
        );

    \I__2381\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11414\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__11431\,
            I => \N__11411\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__11428\,
            I => \N__11408\
        );

    \I__2378\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11401\
        );

    \I__2377\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11401\
        );

    \I__2376\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11401\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__11420\,
            I => d2_count_0
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__11417\,
            I => d2_count_0
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__11414\,
            I => d2_count_0
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__11411\,
            I => d2_count_0
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__11408\,
            I => d2_count_0
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__11401\,
            I => d2_count_0
        );

    \I__2369\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11382\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__11379\,
            I => \N__11376\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__11376\,
            I => \d2.trans_up_1_15\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__11373\,
            I => \d2.trans_up_1_15_cascade_\
        );

    \I__2363\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11367\,
            I => s_dn_0
        );

    \I__2361\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__11361\,
            I => \d1.g2Z0Z_8\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \N__11355\
        );

    \I__2358\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__11352\,
            I => \d1.mins27_0_0\
        );

    \I__2356\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11346\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__11346\,
            I => \d1.g2_i_a5_0Z0Z_7\
        );

    \I__2354\ : InMux
    port map (
            O => \N__11343\,
            I => \N__11339\
        );

    \I__2353\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11336\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11332\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11329\
        );

    \I__2350\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11326\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__11332\,
            I => \N__11323\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__11329\,
            I => d2_trans_up_1_15_1
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__11326\,
            I => d2_trans_up_1_15_1
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__11323\,
            I => d2_trans_up_1_15_1
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__11316\,
            I => \d2_g0_3_cascade_\
        );

    \I__2344\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11310\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__11310\,
            I => \d1.g2_i_a5_1Z0Z_7\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11307\,
            I => \N__11303\
        );

    \I__2341\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11300\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__11303\,
            I => \N__11294\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__11300\,
            I => \N__11294\
        );

    \I__2338\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11291\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__11294\,
            I => \d2.countZ0Z_8\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__11291\,
            I => \d2.countZ0Z_8\
        );

    \I__2335\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11281\
        );

    \I__2334\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11276\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11276\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11273\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11266\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__11273\,
            I => \N__11263\
        );

    \I__2329\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11260\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11255\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11255\
        );

    \I__2326\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11252\
        );

    \I__2325\ : Span4Mux_v
    port map (
            O => \N__11266\,
            I => \N__11249\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__11263\,
            I => d2_trans_up_1_15_8
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__11260\,
            I => d2_trans_up_1_15_8
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__11255\,
            I => d2_trans_up_1_15_8
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__11252\,
            I => d2_trans_up_1_15_8
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__11249\,
            I => d2_trans_up_1_15_8
        );

    \I__2319\ : InMux
    port map (
            O => \N__11238\,
            I => \N__11234\
        );

    \I__2318\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11231\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11225\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11222\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__11230\,
            I => \N__11218\
        );

    \I__2314\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11214\
        );

    \I__2313\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11211\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11208\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__11222\,
            I => \N__11205\
        );

    \I__2310\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11200\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11200\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11197\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__11214\,
            I => \N__11194\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__11211\,
            I => d2_count_6
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__11208\,
            I => d2_count_6
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__11205\,
            I => d2_count_6
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11200\,
            I => d2_count_6
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__11197\,
            I => d2_count_6
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__11194\,
            I => d2_count_6
        );

    \I__2300\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11177\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11174\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__11177\,
            I => \N__11169\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__11174\,
            I => \N__11166\
        );

    \I__2296\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11160\
        );

    \I__2295\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11157\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__11169\,
            I => \N__11154\
        );

    \I__2293\ : Span4Mux_h
    port map (
            O => \N__11166\,
            I => \N__11151\
        );

    \I__2292\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11146\
        );

    \I__2291\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11146\
        );

    \I__2290\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11143\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11140\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__11157\,
            I => d2_count_5
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__11154\,
            I => d2_count_5
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__11151\,
            I => d2_count_5
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__11146\,
            I => d2_count_5
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__11143\,
            I => d2_count_5
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__11140\,
            I => d2_count_5
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__11127\,
            I => \d1.g2_7_0_cascade_\
        );

    \I__2281\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11121\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__11118\,
            I => \d1.g2_11_0\
        );

    \I__2278\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11109\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__11109\,
            I => \d1.N_3\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__11106\,
            I => \N__11103\
        );

    \I__2274\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__11097\,
            I => \N__11094\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__11094\,
            I => \d3.trans_up_1_14_2\
        );

    \I__2270\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11088\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__11085\,
            I => \N__11079\
        );

    \I__2267\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11076\
        );

    \I__2266\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11073\
        );

    \I__2265\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11070\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__11079\,
            I => d3_trans_up_1_15
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__11076\,
            I => d3_trans_up_1_15
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__11073\,
            I => d3_trans_up_1_15
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__11070\,
            I => d3_trans_up_1_15
        );

    \I__2260\ : InMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__11054\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11049\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__11054\,
            I => \N__11046\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11041\
        );

    \I__2255\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11041\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__11049\,
            I => \d1.countZ0Z_5\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__11046\,
            I => \d1.countZ0Z_5\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__11041\,
            I => \d1.countZ0Z_5\
        );

    \I__2251\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__11031\,
            I => \N__11027\
        );

    \I__2249\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11022\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__11027\,
            I => \N__11019\
        );

    \I__2247\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11014\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11014\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__11022\,
            I => \d1.countZ0Z_4\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__11019\,
            I => \d1.countZ0Z_4\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__11014\,
            I => \d1.countZ0Z_4\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__11007\,
            I => \N__11003\
        );

    \I__2241\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10998\
        );

    \I__2240\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10995\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__11002\,
            I => \N__10992\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__11001\,
            I => \N__10989\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10984\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10984\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10979\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10979\
        );

    \I__2233\ : Odrv12
    port map (
            O => \N__10984\,
            I => \d1.countZ0Z_6\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__10979\,
            I => \d1.countZ0Z_6\
        );

    \I__2231\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10970\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10965\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10962\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10957\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10957\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__10965\,
            I => \d1.countZ0Z_3\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__10962\,
            I => \d1.countZ0Z_3\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10957\,
            I => \d1.countZ0Z_3\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10942\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10939\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__10945\,
            I => \N__10936\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__10942\,
            I => \N__10933\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10930\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10927\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__10933\,
            I => \N__10924\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__10930\,
            I => \N__10919\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__10927\,
            I => \N__10919\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__10924\,
            I => \d1.trans_up_1_12\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__10919\,
            I => \d1.trans_up_1_12\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__10914\,
            I => \d1.g1_9_cascade_\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10908\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10908\,
            I => \N__10905\
        );

    \I__2208\ : Odrv12
    port map (
            O => \N__10905\,
            I => \d1.g1_13\
        );

    \I__2207\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10898\
        );

    \I__2206\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10893\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10889\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10886\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10882\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10879\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10875\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__10889\,
            I => \N__10872\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10886\,
            I => \N__10869\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10866\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__10882\,
            I => \N__10861\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__10879\,
            I => \N__10861\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10858\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__10875\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__10872\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__10869\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__10866\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__10861\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10858\,
            I => un1_alarm_on_0_sqmuxa_0
        );

    \I__2188\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10842\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__10842\,
            I => \d1.g2_iZ0Z_0\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__10839\,
            I => \N__10836\
        );

    \I__2185\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10833\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__10833\,
            I => \d1.N_6\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10827\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10827\,
            I => \N__10822\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__10826\,
            I => \N__10819\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10816\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__10822\,
            I => \N__10813\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10810\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__10816\,
            I => ten_secs_1_sqmuxa
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__10813\,
            I => ten_secs_1_sqmuxa
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__10810\,
            I => ten_secs_1_sqmuxa
        );

    \I__2174\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10800\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10800\,
            I => \d1.mins_2_sqmuxa_1\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10794\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__10794\,
            I => \d1.mins_16_1Z0Z_3\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__10791\,
            I => \d1.g3_0_cascade_\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10785\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__10785\,
            I => \d1.N_8_0\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__10782\,
            I => \un1_state_0_sqmuxa_1_0_cascade_\
        );

    \I__2166\ : SRMux
    port map (
            O => \N__10779\,
            I => \N__10775\
        );

    \I__2165\ : CEMux
    port map (
            O => \N__10778\,
            I => \N__10771\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10775\,
            I => \N__10768\
        );

    \I__2163\ : CEMux
    port map (
            O => \N__10774\,
            I => \N__10765\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10771\,
            I => \N__10762\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__10768\,
            I => \N__10759\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__10765\,
            I => \N__10756\
        );

    \I__2159\ : Span4Mux_h
    port map (
            O => \N__10762\,
            I => \N__10753\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__10759\,
            I => \N__10750\
        );

    \I__2157\ : Odrv12
    port map (
            O => \N__10756\,
            I => mins_stored_0_sqmuxa
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__10753\,
            I => mins_stored_0_sqmuxa
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__10750\,
            I => mins_stored_0_sqmuxa
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__10743\,
            I => \N__10740\
        );

    \I__2153\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10737\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10734\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__10734\,
            I => \d1.state_0_sqmuxaZ0Z_1\
        );

    \I__2150\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__10728\,
            I => \N__10725\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__10725\,
            I => \d1.state_0_sqmuxaZ0Z_2\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__10722\,
            I => \d1.state_0_sqmuxaZ0Z_2_cascade_\
        );

    \I__2146\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__10716\,
            I => state_0_sqmuxa
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__10713\,
            I => \state_0_sqmuxa_cascade_\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10706\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10703\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10700\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10697\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__10700\,
            I => \N__10694\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__10697\,
            I => alarm_on_0_sqmuxa
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__10694\,
            I => alarm_on_0_sqmuxa
        );

    \I__2136\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10686\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10683\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__10683\,
            I => \N__10679\
        );

    \I__2133\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10676\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__10679\,
            I => \N__10673\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__10676\,
            I => \alarm_onZ0\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__10673\,
            I => \alarm_onZ0\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10663\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10660\
        );

    \I__2127\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10657\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10663\,
            I => \d3.countZ0Z_16\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10660\,
            I => \d3.countZ0Z_16\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__10657\,
            I => \d3.countZ0Z_16\
        );

    \I__2123\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10645\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10642\
        );

    \I__2121\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10639\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10645\,
            I => \d3.countZ0Z_15\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__10642\,
            I => \d3.countZ0Z_15\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__10639\,
            I => \d3.countZ0Z_15\
        );

    \I__2117\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10627\
        );

    \I__2116\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10624\
        );

    \I__2115\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10621\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__10627\,
            I => \d3.countZ0Z_14\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__10624\,
            I => \d3.countZ0Z_14\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__10621\,
            I => \d3.countZ0Z_14\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10611\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10611\,
            I => \d3.count_RNI4GDSZ0Z_16\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10604\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__10607\,
            I => \N__10601\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10596\
        );

    \I__2106\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10593\
        );

    \I__2105\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10590\
        );

    \I__2104\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10586\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__10596\,
            I => \N__10581\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__10593\,
            I => \N__10581\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__10590\,
            I => \N__10578\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10575\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10572\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__10581\,
            I => \N__10569\
        );

    \I__2097\ : Odrv12
    port map (
            O => \N__10578\,
            I => \ten_secsZ0Z_2\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__10575\,
            I => \ten_secsZ0Z_2\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__10572\,
            I => \ten_secsZ0Z_2\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__10569\,
            I => \ten_secsZ0Z_2\
        );

    \I__2093\ : IoInMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__2091\ : Span4Mux_s3_h
    port map (
            O => \N__10554\,
            I => \N__10551\
        );

    \I__2090\ : Span4Mux_h
    port map (
            O => \N__10551\,
            I => \N__10546\
        );

    \I__2089\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10541\
        );

    \I__2088\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10538\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__10546\,
            I => \N__10535\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__10545\,
            I => \N__10531\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10527\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10541\,
            I => \N__10524\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__10538\,
            I => \N__10519\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__10535\,
            I => \N__10519\
        );

    \I__2081\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10516\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10513\
        );

    \I__2079\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10510\
        );

    \I__2078\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10507\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__10524\,
            I => un1_state_3
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__10519\,
            I => un1_state_3
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10516\,
            I => un1_state_3
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__10513\,
            I => un1_state_3
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10510\,
            I => un1_state_3
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__10507\,
            I => un1_state_3
        );

    \I__2071\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10491\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10491\,
            I => \N__10488\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__10488\,
            I => \N__10485\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__10485\,
            I => \d1.g0_0Z0Z_2\
        );

    \I__2067\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10479\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__10479\,
            I => \N__10475\
        );

    \I__2065\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10470\
        );

    \I__2064\ : Span12Mux_v
    port map (
            O => \N__10475\,
            I => \N__10466\
        );

    \I__2063\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10461\
        );

    \I__2062\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10461\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__10470\,
            I => \N__10458\
        );

    \I__2060\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10455\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__10466\,
            I => \secsZ0Z_2\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__10461\,
            I => \secsZ0Z_2\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__10458\,
            I => \secsZ0Z_2\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__10455\,
            I => \secsZ0Z_2\
        );

    \I__2055\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10437\
        );

    \I__2053\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10432\
        );

    \I__2052\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10427\
        );

    \I__2051\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10427\
        );

    \I__2050\ : Span12Mux_s9_h
    port map (
            O => \N__10437\,
            I => \N__10424\
        );

    \I__2049\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10421\
        );

    \I__2048\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10418\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__10432\,
            I => \secsZ0Z_1\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__10427\,
            I => \secsZ0Z_1\
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__10424\,
            I => \secsZ0Z_1\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__10421\,
            I => \secsZ0Z_1\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__10418\,
            I => \secsZ0Z_1\
        );

    \I__2042\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10404\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__10404\,
            I => \N__10401\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__10401\,
            I => \N__10395\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__10400\,
            I => \N__10392\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__10399\,
            I => \N__10389\
        );

    \I__2037\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10386\
        );

    \I__2036\ : Sp12to4
    port map (
            O => \N__10395\,
            I => \N__10383\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10380\
        );

    \I__2034\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10377\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__10386\,
            I => \secsZ0Z_3\
        );

    \I__2032\ : Odrv12
    port map (
            O => \N__10383\,
            I => \secsZ0Z_3\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__10380\,
            I => \secsZ0Z_3\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__10377\,
            I => \secsZ0Z_3\
        );

    \I__2029\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10365\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__10365\,
            I => \N__10362\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__10362\,
            I => \N__10359\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__10359\,
            I => \N__10353\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10343\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10343\
        );

    \I__2023\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10343\
        );

    \I__2022\ : Span4Mux_h
    port map (
            O => \N__10353\,
            I => \N__10340\
        );

    \I__2021\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10337\
        );

    \I__2020\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10332\
        );

    \I__2019\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10332\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__10343\,
            I => \secsZ0Z_0\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__10340\,
            I => \secsZ0Z_0\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__10337\,
            I => \secsZ0Z_0\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__10332\,
            I => \secsZ0Z_0\
        );

    \I__2014\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10316\
        );

    \I__2012\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10313\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__10316\,
            I => decrement_time_0_secs9
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__10313\,
            I => decrement_time_0_secs9
        );

    \I__2009\ : InMux
    port map (
            O => \N__10308\,
            I => \d2.un3_count_cry_10\
        );

    \I__2008\ : InMux
    port map (
            O => \N__10305\,
            I => \d2.un3_count_cry_11\
        );

    \I__2007\ : InMux
    port map (
            O => \N__10302\,
            I => \d2.un3_count_cry_12\
        );

    \I__2006\ : InMux
    port map (
            O => \N__10299\,
            I => \d2.un3_count_cry_13\
        );

    \I__2005\ : InMux
    port map (
            O => \N__10296\,
            I => \d2.un3_count_cry_14\
        );

    \I__2004\ : InMux
    port map (
            O => \N__10293\,
            I => \d2.un3_count_cry_15\
        );

    \I__2003\ : SRMux
    port map (
            O => \N__10290\,
            I => \N__10281\
        );

    \I__2002\ : SRMux
    port map (
            O => \N__10289\,
            I => \N__10281\
        );

    \I__2001\ : SRMux
    port map (
            O => \N__10288\,
            I => \N__10281\
        );

    \I__2000\ : GlobalMux
    port map (
            O => \N__10281\,
            I => \N__10278\
        );

    \I__1999\ : gio2CtrlBuf
    port map (
            O => \N__10278\,
            I => \d2.idle_i_g\
        );

    \I__1998\ : CEMux
    port map (
            O => \N__10275\,
            I => \N__10272\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10269\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__10269\,
            I => \N__10266\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__10266\,
            I => un1_state_0_sqmuxa_1_0_0
        );

    \I__1994\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10260\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10257\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__10257\,
            I => \d1.state_1_sqmuxaZ0\
        );

    \I__1991\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__10251\,
            I => un1_state_0_sqmuxa_1_0
        );

    \I__1989\ : InMux
    port map (
            O => \N__10248\,
            I => \d2.un3_count_cry_1\
        );

    \I__1988\ : InMux
    port map (
            O => \N__10245\,
            I => \d2.un3_count_cry_2\
        );

    \I__1987\ : InMux
    port map (
            O => \N__10242\,
            I => \d2.un3_count_cry_3\
        );

    \I__1986\ : InMux
    port map (
            O => \N__10239\,
            I => \d2.un3_count_cry_4\
        );

    \I__1985\ : InMux
    port map (
            O => \N__10236\,
            I => \d2.un3_count_cry_5\
        );

    \I__1984\ : InMux
    port map (
            O => \N__10233\,
            I => \d2.un3_count_cry_6\
        );

    \I__1983\ : InMux
    port map (
            O => \N__10230\,
            I => \d2.un3_count_cry_7\
        );

    \I__1982\ : InMux
    port map (
            O => \N__10227\,
            I => \bfn_11_19_0_\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10224\,
            I => \d2.un3_count_cry_9\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__10218\,
            I => \N__10214\
        );

    \I__1978\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__1977\ : Odrv12
    port map (
            O => \N__10214\,
            I => \d1.trans_up_1_0\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__10211\,
            I => \d1.trans_up_1_0\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__1974\ : InMux
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__10200\,
            I => \d1.g2_i_a5_3\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__10197\,
            I => \d1.g0_0_0Z0Z_1_cascade_\
        );

    \I__1971\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10191\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__10191\,
            I => \d1.g2Z0Z_10\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__10188\,
            I => \N__10184\
        );

    \I__1968\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10181\
        );

    \I__1967\ : InMux
    port map (
            O => \N__10184\,
            I => \N__10178\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__10181\,
            I => \N__10175\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10172\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__10175\,
            I => \d1.g0_2_0_a4Z0Z_2\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__10172\,
            I => \d1.g0_2_0_a4Z0Z_2\
        );

    \I__1962\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10164\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__10164\,
            I => \N__10158\
        );

    \I__1960\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10155\
        );

    \I__1959\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10150\
        );

    \I__1958\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10147\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__10158\,
            I => \N__10144\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__10155\,
            I => \N__10141\
        );

    \I__1955\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10136\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10136\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__10150\,
            I => s_dn
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__10147\,
            I => s_dn
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__10144\,
            I => s_dn
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__10141\,
            I => s_dn
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10136\,
            I => s_dn
        );

    \I__1948\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10121\
        );

    \I__1947\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10118\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__10121\,
            I => \d1.g0_2_0_o2_2\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__10118\,
            I => \d1.g0_2_0_o2_2\
        );

    \I__1944\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10110\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10107\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__10107\,
            I => \d1.g2_i_a5_0Z0Z_3\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__10104\,
            I => \d1.g2_i_a5_0Z0Z_6_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10098\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__10098\,
            I => \d1.g2_i_a5Z0Z_2\
        );

    \I__1938\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__10089\,
            I => \d1.secs_0_sqmuxa_xZ0Z1\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__1934\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10080\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10077\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__10077\,
            I => \N__10074\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__10074\,
            I => \N__10071\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__10071\,
            I => \mins_storedZ0Z_3\
        );

    \I__1929\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10065\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10065\,
            I => \d1.N_5\
        );

    \I__1927\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10056\
        );

    \I__1926\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10053\
        );

    \I__1925\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10048\
        );

    \I__1924\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10048\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__10056\,
            I => \d1.un1_mins_1_sqmuxa_0\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__10053\,
            I => \d1.un1_mins_1_sqmuxa_0\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__10048\,
            I => \d1.un1_mins_1_sqmuxa_0\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10038\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__10035\,
            I => \d1.g0_0_0_a4_2_1\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__10032\,
            I => \secs_RNO_0Z0Z_2_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10026\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__10026\,
            I => \N__10020\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10017\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10014\
        );

    \I__1912\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10011\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__10020\,
            I => secs_0_sqmuxa
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__10017\,
            I => secs_0_sqmuxa
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__10014\,
            I => secs_0_sqmuxa
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__10011\,
            I => secs_0_sqmuxa
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__10002\,
            I => \N__9996\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__10001\,
            I => \N__9993\
        );

    \I__1905\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9984\
        );

    \I__1904\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9984\
        );

    \I__1903\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9984\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9984\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9984\,
            I => un1_state_7_0
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__9981\,
            I => \un1_secs_c3_cascade_\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9969\
        );

    \I__1898\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9969\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9969\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9969\,
            I => un1_alarm_on_0_sqmuxa_0_i
        );

    \I__1895\ : InMux
    port map (
            O => \N__9966\,
            I => \d3.un3_count_cry_14\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9963\,
            I => \d3.un3_count_cry_15\
        );

    \I__1893\ : SRMux
    port map (
            O => \N__9960\,
            I => \N__9951\
        );

    \I__1892\ : SRMux
    port map (
            O => \N__9959\,
            I => \N__9951\
        );

    \I__1891\ : SRMux
    port map (
            O => \N__9958\,
            I => \N__9951\
        );

    \I__1890\ : GlobalMux
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__1889\ : gio2CtrlBuf
    port map (
            O => \N__9948\,
            I => \d3.idle_i_g\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9935\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9920\
        );

    \I__1886\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9920\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9920\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9920\
        );

    \I__1883\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9920\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9920\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9920\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__9935\,
            I => \N__9912\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9908\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9897\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9897\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9897\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9897\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9897\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__9912\,
            I => \N__9894\
        );

    \I__1872\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9891\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__9908\,
            I => \decrement_time_0_prescaler10_THRU_CO\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9897\,
            I => \decrement_time_0_prescaler10_THRU_CO\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__9894\,
            I => \decrement_time_0_prescaler10_THRU_CO\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__9891\,
            I => \decrement_time_0_prescaler10_THRU_CO\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__9882\,
            I => \un1_state_7_0_cascade_\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__9879\,
            I => \un1_alarm_on_0_sqmuxa_0_i_cascade_\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9876\,
            I => \N__9873\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N_120_1\
        );

    \I__1863\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9862\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9859\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9854\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9854\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9851\
        );

    \I__1858\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9848\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__9862\,
            I => s_cancel
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__9859\,
            I => s_cancel
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__9854\,
            I => s_cancel
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__9851\,
            I => s_cancel
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__9848\,
            I => s_cancel
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__9837\,
            I => \N__9833\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9829\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9826\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9823\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9829\,
            I => \d3.countZ0Z_13\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__9826\,
            I => \d3.countZ0Z_13\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__9823\,
            I => \d3.countZ0Z_13\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9813\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9813\,
            I => \N__9809\
        );

    \I__1843\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9806\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__9809\,
            I => d3_g0_1
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__9806\,
            I => d3_g0_1
        );

    \I__1840\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9797\
        );

    \I__1839\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9794\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__9797\,
            I => \d3.countZ0Z_6\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__9794\,
            I => \d3.countZ0Z_6\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9789\,
            I => \d3.un3_count_cry_5\
        );

    \I__1835\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9782\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9779\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__9782\,
            I => \d3.countZ0Z_7\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__9779\,
            I => \d3.countZ0Z_7\
        );

    \I__1831\ : InMux
    port map (
            O => \N__9774\,
            I => \d3.un3_count_cry_6\
        );

    \I__1830\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9767\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9764\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__9767\,
            I => \d3.countZ0Z_8\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__9764\,
            I => \d3.countZ0Z_8\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9759\,
            I => \d3.un3_count_cry_7\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__9756\,
            I => \N__9752\
        );

    \I__1824\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9749\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9746\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__9749\,
            I => \d3.countZ0Z_9\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__9746\,
            I => \d3.countZ0Z_9\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9741\,
            I => \bfn_11_14_0_\
        );

    \I__1819\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9734\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9731\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9728\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__9731\,
            I => \d3.countZ0Z_10\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__9728\,
            I => \d3.countZ0Z_10\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9723\,
            I => \d3.un3_count_cry_9\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__9720\,
            I => \N__9717\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9713\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9710\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__9713\,
            I => \N__9707\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9710\,
            I => \d3.countZ0Z_11\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__9707\,
            I => \d3.countZ0Z_11\
        );

    \I__1807\ : InMux
    port map (
            O => \N__9702\,
            I => \d3.un3_count_cry_10\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__9699\,
            I => \N__9696\
        );

    \I__1805\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9692\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9689\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__9692\,
            I => \N__9686\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__9689\,
            I => \d3.countZ0Z_12\
        );

    \I__1801\ : Odrv12
    port map (
            O => \N__9686\,
            I => \d3.countZ0Z_12\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9681\,
            I => \d3.un3_count_cry_11\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9678\,
            I => \d3.un3_count_cry_12\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9675\,
            I => \d3.un3_count_cry_13\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__9672\,
            I => \N__9668\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9665\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9662\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__9665\,
            I => \d4.countZ0Z_14\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__9662\,
            I => \d4.countZ0Z_14\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9657\,
            I => \d4.un3_count_cry_13\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9650\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9647\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__9650\,
            I => \d4.countZ0Z_15\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__9647\,
            I => \d4.countZ0Z_15\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9642\,
            I => \d4.un3_count_cry_14\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9639\,
            I => \d4.un3_count_cry_15\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__9636\,
            I => \N__9632\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9629\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9626\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__9629\,
            I => \d4.countZ0Z_16\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__9626\,
            I => \d4.countZ0Z_16\
        );

    \I__1780\ : SRMux
    port map (
            O => \N__9621\,
            I => \N__9612\
        );

    \I__1779\ : SRMux
    port map (
            O => \N__9620\,
            I => \N__9612\
        );

    \I__1778\ : SRMux
    port map (
            O => \N__9619\,
            I => \N__9612\
        );

    \I__1777\ : GlobalMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__1776\ : gio2CtrlBuf
    port map (
            O => \N__9609\,
            I => \d4.idle_i_g\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9600\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9593\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9593\
        );

    \I__1772\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9593\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__9600\,
            I => \d3.countZ0Z_0\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__9593\,
            I => \d3.countZ0Z_0\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__9588\,
            I => \N__9584\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__9587\,
            I => \N__9581\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9577\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9572\
        );

    \I__1765\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9572\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__9577\,
            I => \d3.countZ0Z_1\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__9572\,
            I => \d3.countZ0Z_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9563\
        );

    \I__1761\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__9563\,
            I => \d3.countZ0Z_2\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__9560\,
            I => \d3.countZ0Z_2\
        );

    \I__1758\ : InMux
    port map (
            O => \N__9555\,
            I => \d3.un3_count_cry_1\
        );

    \I__1757\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9548\
        );

    \I__1756\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9545\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9548\,
            I => \d3.countZ0Z_3\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__9545\,
            I => \d3.countZ0Z_3\
        );

    \I__1753\ : InMux
    port map (
            O => \N__9540\,
            I => \d3.un3_count_cry_2\
        );

    \I__1752\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9533\
        );

    \I__1751\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9530\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__9533\,
            I => \d3.countZ0Z_4\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__9530\,
            I => \d3.countZ0Z_4\
        );

    \I__1748\ : InMux
    port map (
            O => \N__9525\,
            I => \d3.un3_count_cry_3\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__9522\,
            I => \N__9518\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9515\
        );

    \I__1745\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9512\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__9515\,
            I => \d3.countZ0Z_5\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__9512\,
            I => \d3.countZ0Z_5\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9507\,
            I => \d3.un3_count_cry_4\
        );

    \I__1741\ : InMux
    port map (
            O => \N__9504\,
            I => \d4.un3_count_cry_4\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__9501\,
            I => \N__9497\
        );

    \I__1739\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9494\
        );

    \I__1738\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9491\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__9494\,
            I => \d4.countZ0Z_6\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__9491\,
            I => \d4.countZ0Z_6\
        );

    \I__1735\ : InMux
    port map (
            O => \N__9486\,
            I => \d4.un3_count_cry_5\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9479\
        );

    \I__1733\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9476\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__9479\,
            I => \d4.countZ0Z_7\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__9476\,
            I => \d4.countZ0Z_7\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9471\,
            I => \d4.un3_count_cry_6\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9464\
        );

    \I__1728\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9461\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__9464\,
            I => \d4.countZ0Z_8\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__9461\,
            I => \d4.countZ0Z_8\
        );

    \I__1725\ : InMux
    port map (
            O => \N__9456\,
            I => \d4.un3_count_cry_7\
        );

    \I__1724\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9449\
        );

    \I__1723\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9446\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__9449\,
            I => \d4.countZ0Z_9\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__9446\,
            I => \d4.countZ0Z_9\
        );

    \I__1720\ : InMux
    port map (
            O => \N__9441\,
            I => \bfn_11_12_0_\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__9438\,
            I => \N__9434\
        );

    \I__1718\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9431\
        );

    \I__1717\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9428\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__9431\,
            I => \d4.countZ0Z_10\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__9428\,
            I => \d4.countZ0Z_10\
        );

    \I__1714\ : InMux
    port map (
            O => \N__9423\,
            I => \d4.un3_count_cry_9\
        );

    \I__1713\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9416\
        );

    \I__1712\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9413\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9416\,
            I => \d4.countZ0Z_11\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__9413\,
            I => \d4.countZ0Z_11\
        );

    \I__1709\ : InMux
    port map (
            O => \N__9408\,
            I => \d4.un3_count_cry_10\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__9405\,
            I => \N__9401\
        );

    \I__1707\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9398\
        );

    \I__1706\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9395\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__9398\,
            I => \d4.countZ0Z_12\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__9395\,
            I => \d4.countZ0Z_12\
        );

    \I__1703\ : InMux
    port map (
            O => \N__9390\,
            I => \d4.un3_count_cry_11\
        );

    \I__1702\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9383\
        );

    \I__1701\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9380\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__9383\,
            I => \d4.countZ0Z_13\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__9380\,
            I => \d4.countZ0Z_13\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9375\,
            I => \d4.un3_count_cry_12\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__9372\,
            I => \d1.g2Z0Z_7_cascade_\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__9369\,
            I => \d1.g0_1_0_a4Z0Z_7_cascade_\
        );

    \I__1695\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9363\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__9363\,
            I => \N__9357\
        );

    \I__1693\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9352\
        );

    \I__1692\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9352\
        );

    \I__1691\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9349\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__9357\,
            I => \N__9346\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__9352\,
            I => \d4.countZ0Z_0\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__9349\,
            I => \d4.countZ0Z_0\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__9346\,
            I => \d4.countZ0Z_0\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__9339\,
            I => \N__9334\
        );

    \I__1685\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9331\
        );

    \I__1684\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9328\
        );

    \I__1683\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9325\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9322\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__9328\,
            I => \d4.countZ0Z_1\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__9325\,
            I => \d4.countZ0Z_1\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__9322\,
            I => \d4.countZ0Z_1\
        );

    \I__1678\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9311\
        );

    \I__1677\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9308\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__9311\,
            I => \d4.countZ0Z_2\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9308\,
            I => \d4.countZ0Z_2\
        );

    \I__1674\ : InMux
    port map (
            O => \N__9303\,
            I => \d4.un3_count_cry_1\
        );

    \I__1673\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9296\
        );

    \I__1672\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9293\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__9296\,
            I => \d4.countZ0Z_3\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__9293\,
            I => \d4.countZ0Z_3\
        );

    \I__1669\ : InMux
    port map (
            O => \N__9288\,
            I => \d4.un3_count_cry_2\
        );

    \I__1668\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9281\
        );

    \I__1667\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9278\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__9281\,
            I => \d4.countZ0Z_4\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__9278\,
            I => \d4.countZ0Z_4\
        );

    \I__1664\ : InMux
    port map (
            O => \N__9273\,
            I => \d4.un3_count_cry_3\
        );

    \I__1663\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9266\
        );

    \I__1662\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9263\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__9266\,
            I => \d4.countZ0Z_5\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__9263\,
            I => \d4.countZ0Z_5\
        );

    \I__1659\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__9255\,
            I => \N__9252\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__9252\,
            I => \d1.g2_8_1\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__9249\,
            I => \d2.g0_0_10_cascade_\
        );

    \I__1655\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__9243\,
            I => \d2.g0_0_12\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \d2.g0_0_14_cascade_\
        );

    \I__1652\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__9231\,
            I => \d1.g2_8_0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__9225\,
            I => \d2.g0_0_11\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__1646\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__9216\,
            I => \d2.trans_up_1_14_2\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9210\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__9210\,
            I => \d1.g1_7\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__1641\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__9201\,
            I => \d1.g1_8\
        );

    \I__1639\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__9195\,
            I => \d1.g1_14\
        );

    \I__1637\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__9183\,
            I => \d1.g0_1_a5_0_10\
        );

    \I__1633\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__9174\,
            I => \d1.g0_1_a5_0_15\
        );

    \I__1630\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9164\
        );

    \I__1628\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9161\
        );

    \I__1627\ : Span4Mux_h
    port map (
            O => \N__9164\,
            I => \N__9158\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__9161\,
            I => \d1.trans_up_1_10\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__9158\,
            I => \d1.trans_up_1_10\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__9153\,
            I => \N__9149\
        );

    \I__1623\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9146\
        );

    \I__1622\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__9146\,
            I => \N__9140\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__9143\,
            I => \N__9137\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__9140\,
            I => \N__9132\
        );

    \I__1618\ : Span4Mux_h
    port map (
            O => \N__9137\,
            I => \N__9132\
        );

    \I__1617\ : Span4Mux_h
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__9129\,
            I => \d1.trans_up_1_11\
        );

    \I__1615\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__9120\,
            I => \N__9116\
        );

    \I__1612\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9113\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__9116\,
            I => \d1.trans_up_1_13\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__9113\,
            I => \d1.trans_up_1_13\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__9108\,
            I => \d1.trans_up_1_0_cascade_\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__9105\,
            I => \d1.g0_2_0_o2_2_cascade_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__9099\,
            I => \N__9096\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__9093\,
            I => \mins_storedZ0Z_0\
        );

    \I__1603\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__9087\,
            I => \d1.g0_0_0\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__9084\,
            I => \d1.N_19_i_cascade_\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__9081\,
            I => \N__9077\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9073\
        );

    \I__1598\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9070\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__9076\,
            I => \N__9067\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9060\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9060\
        );

    \I__1594\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9057\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__9066\,
            I => \N__9053\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9049\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__9060\,
            I => \N__9043\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9043\
        );

    \I__1589\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9038\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9038\
        );

    \I__1587\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9035\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9049\,
            I => \N__9032\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9029\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__9043\,
            I => \N__9026\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__9038\,
            I => \N__9023\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__9035\,
            I => \d1.stateZ0Z_0\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__9032\,
            I => \d1.stateZ0Z_0\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__9029\,
            I => \d1.stateZ0Z_0\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__9026\,
            I => \d1.stateZ0Z_0\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__9023\,
            I => \d1.stateZ0Z_0\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__9012\,
            I => \N__9009\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__1574\ : Odrv12
    port map (
            O => \N__9003\,
            I => \d1.ten_secs_1_sqmuxa_0\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8997\,
            I => \d1.g2_0Z0Z_4\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8991\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8988\
        );

    \I__1569\ : Odrv12
    port map (
            O => \N__8988\,
            I => \d1.g2_0Z0Z_3\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__8985\,
            I => \ten_secs_1_sqmuxa_cascade_\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8979\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__1565\ : Odrv12
    port map (
            O => \N__8976\,
            I => \d1.g1_0\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__8973\,
            I => \d1.g0_0_0_0_0_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__8967\,
            I => \mins_storedZ0Z_1\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__8964\,
            I => \d1.un1_mins_4_0_1_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8957\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8953\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8950\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8947\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8944\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__8950\,
            I => \N__8941\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__8947\,
            I => \d1.countZ0Z_9\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__8944\,
            I => \d1.countZ0Z_9\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__8941\,
            I => \d1.countZ0Z_9\
        );

    \I__1551\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8930\
        );

    \I__1550\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8926\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8923\
        );

    \I__1548\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8920\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__8926\,
            I => \N__8917\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__8923\,
            I => \N__8914\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__8920\,
            I => \d1.countZ0Z_8\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__8917\,
            I => \d1.countZ0Z_8\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__8914\,
            I => \d1.countZ0Z_8\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8900\
        );

    \I__1540\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8896\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8893\
        );

    \I__1538\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8890\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__8896\,
            I => \N__8887\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__8893\,
            I => \N__8884\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__8890\,
            I => \d1.countZ0Z_10\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__8887\,
            I => \d1.countZ0Z_10\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__8884\,
            I => \d1.countZ0Z_10\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8872\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8869\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8866\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__8872\,
            I => \N__8863\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8869\,
            I => \N__8858\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__8866\,
            I => \N__8858\
        );

    \I__1526\ : Span4Mux_h
    port map (
            O => \N__8863\,
            I => \N__8855\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__8858\,
            I => \d1.countZ0Z_7\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__8855\,
            I => \d1.countZ0Z_7\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8846\
        );

    \I__1522\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8843\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__8846\,
            I => \d1.trans_up_1_9\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8843\,
            I => \d1.trans_up_1_9\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8835\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8835\,
            I => \d1.g2Z0Z_11\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__8832\,
            I => \d1.un1_mins_1_sqmuxa_0_cascade_\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__8829\,
            I => \d1.un1_mins_3_sqmuxa_0_0_cascade_\
        );

    \I__1515\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__8823\,
            I => \d1.N_4\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8817\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8814\
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__8814\,
            I => \mins_storedZ0Z_2\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__8811\,
            I => \d1.g1_cascade_\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__8808\,
            I => \d4_trans_up_1_cascade_\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__8805\,
            I => \ten_secs_r_1_1_cascade_\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__8802\,
            I => \d3.trans_up_1_14_2_cascade_\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__8799\,
            I => \s_cancel_cascade_\
        );

    \I__1505\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8789\
        );

    \I__1504\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8786\
        );

    \I__1503\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8779\
        );

    \I__1502\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8779\
        );

    \I__1501\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8779\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8776\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8773\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__8779\,
            I => \N__8770\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__8776\,
            I => d4_state
        );

    \I__1496\ : Odrv12
    port map (
            O => \N__8773\,
            I => d4_state
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__8770\,
            I => d4_state
        );

    \I__1494\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8759\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8756\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__8759\,
            I => d4_trans_up_1
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__8756\,
            I => d4_trans_up_1
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__8751\,
            I => \secs_0_sqmuxa_cascade_\
        );

    \I__1489\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8744\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8740\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8737\
        );

    \I__1486\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8734\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__8740\,
            I => un1_state_9_0
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__8737\,
            I => un1_state_9_0
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__8734\,
            I => un1_state_9_0
        );

    \I__1482\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__8724\,
            I => \d3.trans_up_1_15_8\
        );

    \I__1480\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8717\
        );

    \I__1479\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8714\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8709\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8709\
        );

    \I__1476\ : Odrv12
    port map (
            O => \N__8709\,
            I => \d4.syncZ0Z_1\
        );

    \I__1475\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__8703\,
            I => \d3.trans_up_1_15_7\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8694\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__8694\,
            I => \d4.trans_up_1_9\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__8688\,
            I => \d4.trans_up_1_12\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__8682\,
            I => \d4.trans_up_1_11\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__8679\,
            I => \d4.trans_up_1_13_cascade_\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__8673\,
            I => \d4.trans_up_1_10\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__8670\,
            I => \d1.g2Z0Z_1_cascade_\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__8667\,
            I => \d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8659\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8656\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8652\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__8659\,
            I => \N__8649\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8646\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8643\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8652\,
            I => \N__8640\
        );

    \I__1454\ : Span4Mux_v
    port map (
            O => \N__8649\,
            I => \N__8635\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8635\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__8643\,
            I => \a.countZ0Z_0\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__8640\,
            I => \a.countZ0Z_0\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__8635\,
            I => \a.countZ0Z_0\
        );

    \I__1449\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__8622\,
            I => \d3.trans_up_1_15_1\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1445\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8607\
        );

    \I__1443\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8604\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8601\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8598\
        );

    \I__1440\ : Span4Mux_h
    port map (
            O => \N__8607\,
            I => \N__8595\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8592\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8589\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__8598\,
            I => \d1.countZ0Z_12\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__8595\,
            I => \d1.countZ0Z_12\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__8592\,
            I => \d1.countZ0Z_12\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__8589\,
            I => \d1.countZ0Z_12\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8577\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1430\ : Sp12to4
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__1429\ : Span12Mux_h
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1428\ : Odrv12
    port map (
            O => \N__8565\,
            I => switch_cancel_c
        );

    \I__1427\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__8553\,
            I => \d3.syncZ0Z_0\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1421\ : Odrv12
    port map (
            O => \N__8544\,
            I => \d1.g2_7_1\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__8532\,
            I => \d2.syncZ0Z_0\
        );

    \I__1416\ : IoInMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__1414\ : IoSpan4Mux
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1413\ : Span4Mux_s2_v
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__8511\,
            I => \d4.idle_i\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__8505\,
            I => \d1.g2_12_0\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__8502\,
            I => \d1.g2Z0Z_12_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8492\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8489\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__8492\,
            I => \N__8486\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__8489\,
            I => \prescalerZ0Z_10\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__8486\,
            I => \prescalerZ0Z_10\
        );

    \I__1400\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8477\
        );

    \I__1399\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8474\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__8477\,
            I => \prescalerZ0Z_11\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__8474\,
            I => \prescalerZ0Z_11\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__8469\,
            I => \N__8465\
        );

    \I__1395\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8462\
        );

    \I__1394\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8459\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__8462\,
            I => \prescalerZ0Z_9\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__8459\,
            I => \prescalerZ0Z_9\
        );

    \I__1391\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8450\
        );

    \I__1390\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8447\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__8450\,
            I => \prescalerZ0Z_12\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__8447\,
            I => \prescalerZ0Z_12\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__8442\,
            I => \N__8439\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__8430\,
            I => decrement_time_0_prescaler10_5_and
        );

    \I__1382\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8423\
        );

    \I__1381\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8420\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__8423\,
            I => \N__8417\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__8420\,
            I => \prescalerZ0Z_25\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__8417\,
            I => \prescalerZ0Z_25\
        );

    \I__1377\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8408\
        );

    \I__1376\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8405\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__8408\,
            I => \prescalerZ0Z_27\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8405\,
            I => \prescalerZ0Z_27\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__8400\,
            I => \N__8396\
        );

    \I__1372\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8393\
        );

    \I__1371\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8390\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__8393\,
            I => \prescalerZ0Z_17\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__8390\,
            I => \prescalerZ0Z_17\
        );

    \I__1368\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8381\
        );

    \I__1367\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8378\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__8381\,
            I => \prescalerZ0Z_19\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__8378\,
            I => \prescalerZ0Z_19\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__1363\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__8361\,
            I => decrement_time_0_prescaler10_6_and
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__8358\,
            I => \d1.g2_7_2_cascade_\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__8355\,
            I => \d1.mins27_1_cascade_\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__8352\,
            I => \d1.g2Z0Z_0_cascade_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__8346\,
            I => \N__8343\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__8343\,
            I => \d1.g0_1_a5_0_9\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8337\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__8334\,
            I => \d1.g0_1_a5_0_8\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__8325\,
            I => \d1.g0_0_0_a4_2_0\
        );

    \I__1347\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__8319\,
            I => \d1.gZ0Z2\
        );

    \I__1345\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8310\
        );

    \I__1344\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8310\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8305\
        );

    \I__1342\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8300\
        );

    \I__1341\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8297\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__8305\,
            I => \N__8294\
        );

    \I__1339\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8289\
        );

    \I__1338\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8289\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__8300\,
            I => \d1.countZ0Z_0\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__8297\,
            I => \d1.countZ0Z_0\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__8294\,
            I => \d1.countZ0Z_0\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__8289\,
            I => \d1.countZ0Z_0\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__1332\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8271\
        );

    \I__1331\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8271\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__8271\,
            I => \N__8266\
        );

    \I__1329\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8263\
        );

    \I__1328\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8260\
        );

    \I__1327\ : Span4Mux_h
    port map (
            O => \N__8266\,
            I => \N__8257\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__8263\,
            I => \N__8254\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__8260\,
            I => \d1.countZ0Z_11\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__8257\,
            I => \d1.countZ0Z_11\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__8254\,
            I => \d1.countZ0Z_11\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1321\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__8241\,
            I => decrement_time_0_prescaler10_2_and
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1318\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__8232\,
            I => decrement_time_0_prescaler10_3_and
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__1315\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__8220\,
            I => decrement_time_0_prescaler10_4_and
        );

    \I__1312\ : InMux
    port map (
            O => \N__8217\,
            I => decrement_time_0_prescaler10
        );

    \I__1311\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1309\ : Span4Mux_h
    port map (
            O => \N__8208\,
            I => \N__8205\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__8205\,
            I => \prescaler_1_cry_12_THRU_CO\
        );

    \I__1307\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8194\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8191\
        );

    \I__1304\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8188\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__8194\,
            I => \N__8185\
        );

    \I__1302\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8182\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__8188\,
            I => \prescalerZ0Z_13\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__8185\,
            I => \prescalerZ0Z_13\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__8182\,
            I => \prescalerZ0Z_13\
        );

    \I__1298\ : InMux
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__8166\,
            I => \prescaler_1_cry_13_THRU_CO\
        );

    \I__1294\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__8157\,
            I => \N__8152\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8147\
        );

    \I__1290\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8147\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__8152\,
            I => \prescalerZ0Z_14\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__8147\,
            I => \prescalerZ0Z_14\
        );

    \I__1287\ : InMux
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__8130\,
            I => \prescaler_1_cry_14_THRU_CO\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__8121\,
            I => \N__8116\
        );

    \I__1279\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8111\
        );

    \I__1278\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8111\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__8116\,
            I => \prescalerZ0Z_15\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__8111\,
            I => \prescalerZ0Z_15\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__8097\,
            I => \prescaler_1_cry_15_THRU_CO\
        );

    \I__1271\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__8091\,
            I => \N__8087\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__8090\,
            I => \N__8084\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__8087\,
            I => \N__8080\
        );

    \I__1267\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8075\
        );

    \I__1266\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8075\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__8080\,
            I => \prescalerZ0Z_16\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8075\,
            I => \prescalerZ0Z_16\
        );

    \I__1263\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__8061\,
            I => \prescaler_1_cry_17_THRU_CO\
        );

    \I__1259\ : CEMux
    port map (
            O => \N__8058\,
            I => \N__8037\
        );

    \I__1258\ : CEMux
    port map (
            O => \N__8057\,
            I => \N__8037\
        );

    \I__1257\ : CEMux
    port map (
            O => \N__8056\,
            I => \N__8037\
        );

    \I__1256\ : CEMux
    port map (
            O => \N__8055\,
            I => \N__8037\
        );

    \I__1255\ : CEMux
    port map (
            O => \N__8054\,
            I => \N__8037\
        );

    \I__1254\ : CEMux
    port map (
            O => \N__8053\,
            I => \N__8037\
        );

    \I__1253\ : CEMux
    port map (
            O => \N__8052\,
            I => \N__8037\
        );

    \I__1252\ : GlobalMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1251\ : gio2CtrlBuf
    port map (
            O => \N__8034\,
            I => un1_state_3_g
        );

    \I__1250\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8024\
        );

    \I__1248\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8020\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__8024\,
            I => \N__8017\
        );

    \I__1246\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8014\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__8020\,
            I => \prescalerZ0Z_20\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__8017\,
            I => \prescalerZ0Z_20\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__8014\,
            I => \prescalerZ0Z_20\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__8000\
        );

    \I__1240\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7996\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__8000\,
            I => \N__7993\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7990\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__7996\,
            I => \prescalerZ0Z_21\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__7993\,
            I => \prescalerZ0Z_21\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7990\,
            I => \prescalerZ0Z_21\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7976\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__7979\,
            I => \N__7973\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7969\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7966\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7963\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__7969\,
            I => \N__7958\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__7966\,
            I => \N__7958\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7963\,
            I => \prescalerZ0Z_22\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__7958\,
            I => \prescalerZ0Z_22\
        );

    \I__1224\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__7947\,
            I => \N__7942\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7937\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7937\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__7942\,
            I => \prescalerZ0Z_18\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7937\,
            I => \prescalerZ0Z_18\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1216\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__7926\,
            I => decrement_time_0_prescaler10_0_and
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__7917\,
            I => decrement_time_0_prescaler10_1_and
        );

    \I__1211\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__7911\,
            I => \N__7908\
        );

    \I__1209\ : Span12Mux_v
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__7905\,
            I => \prescaler_1_cry_7_THRU_CO\
        );

    \I__1207\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7898\
        );

    \I__1206\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7895\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7892\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7895\,
            I => \N__7886\
        );

    \I__1203\ : Span4Mux_v
    port map (
            O => \N__7892\,
            I => \N__7886\
        );

    \I__1202\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7883\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__7886\,
            I => \prescalerZ0Z_8\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__7883\,
            I => \prescalerZ0Z_8\
        );

    \I__1199\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__7869\,
            I => \prescaler_1_cry_22_THRU_CO\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__7860\,
            I => \N__7855\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7850\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7850\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__7855\,
            I => \prescalerZ0Z_23\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7850\,
            I => \prescalerZ0Z_23\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__7836\,
            I => \prescaler_1_cry_23_THRU_CO\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7825\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__7829\,
            I => \N__7822\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7819\
        );

    \I__1180\ : Sp12to4
    port map (
            O => \N__7825\,
            I => \N__7816\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7813\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__7819\,
            I => \prescalerZ0Z_24\
        );

    \I__1177\ : Odrv12
    port map (
            O => \N__7816\,
            I => \prescalerZ0Z_24\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7813\,
            I => \prescalerZ0Z_24\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1173\ : Span4Mux_h
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__7794\,
            I => \prescaler_1_cry_25_THRU_CO\
        );

    \I__1170\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__7788\,
            I => \N__7785\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__7785\,
            I => \N__7780\
        );

    \I__1167\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7775\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7775\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__7780\,
            I => \prescalerZ0Z_26\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7775\,
            I => \prescalerZ0Z_26\
        );

    \I__1163\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__7758\,
            I => \prescaler_1_cry_19_THRU_CO\
        );

    \I__1158\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7752\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__7749\,
            I => \N__7746\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__7746\,
            I => \prescaler_1_cry_20_THRU_CO\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7737\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__7734\,
            I => \prescaler_1_cry_21_THRU_CO\
        );

    \I__1150\ : InMux
    port map (
            O => \N__7731\,
            I => prescaler_1_cry_18
        );

    \I__1149\ : InMux
    port map (
            O => \N__7728\,
            I => prescaler_1_cry_19
        );

    \I__1148\ : InMux
    port map (
            O => \N__7725\,
            I => prescaler_1_cry_20
        );

    \I__1147\ : InMux
    port map (
            O => \N__7722\,
            I => prescaler_1_cry_21
        );

    \I__1146\ : InMux
    port map (
            O => \N__7719\,
            I => prescaler_1_cry_22
        );

    \I__1145\ : InMux
    port map (
            O => \N__7716\,
            I => prescaler_1_cry_23
        );

    \I__1144\ : InMux
    port map (
            O => \N__7713\,
            I => \bfn_8_18_0_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7710\,
            I => prescaler_1_cry_25
        );

    \I__1142\ : InMux
    port map (
            O => \N__7707\,
            I => prescaler_1_cry_26
        );

    \I__1141\ : InMux
    port map (
            O => \N__7704\,
            I => prescaler_1_cry_9
        );

    \I__1140\ : InMux
    port map (
            O => \N__7701\,
            I => prescaler_1_cry_10
        );

    \I__1139\ : InMux
    port map (
            O => \N__7698\,
            I => prescaler_1_cry_11
        );

    \I__1138\ : InMux
    port map (
            O => \N__7695\,
            I => prescaler_1_cry_12
        );

    \I__1137\ : InMux
    port map (
            O => \N__7692\,
            I => prescaler_1_cry_13
        );

    \I__1136\ : InMux
    port map (
            O => \N__7689\,
            I => prescaler_1_cry_14
        );

    \I__1135\ : InMux
    port map (
            O => \N__7686\,
            I => prescaler_1_cry_15
        );

    \I__1134\ : InMux
    port map (
            O => \N__7683\,
            I => \bfn_8_17_0_\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7680\,
            I => prescaler_1_cry_17
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__7677\,
            I => \N__7671\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7666\
        );

    \I__1130\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7666\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7663\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7671\,
            I => \N__7660\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7666\,
            I => \prescalerZ0Z_0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__7663\,
            I => \prescalerZ0Z_0\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__7660\,
            I => \prescalerZ0Z_0\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__7653\,
            I => \N__7649\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7645\
        );

    \I__1122\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7642\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7648\,
            I => \N__7639\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7645\,
            I => \prescalerZ0Z_1\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7642\,
            I => \prescalerZ0Z_1\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__7639\,
            I => \prescalerZ0Z_1\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7628\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7631\,
            I => \N__7625\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7622\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7625\,
            I => \prescalerZ0Z_2\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__7622\,
            I => \prescalerZ0Z_2\
        );

    \I__1112\ : InMux
    port map (
            O => \N__7617\,
            I => prescaler_1_cry_1
        );

    \I__1111\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7610\
        );

    \I__1110\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7607\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__7610\,
            I => \N__7604\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__7607\,
            I => \prescalerZ0Z_3\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__7604\,
            I => \prescalerZ0Z_3\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7599\,
            I => prescaler_1_cry_2
        );

    \I__1105\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7592\
        );

    \I__1104\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7589\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7592\,
            I => \prescalerZ0Z_4\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__7589\,
            I => \prescalerZ0Z_4\
        );

    \I__1101\ : InMux
    port map (
            O => \N__7584\,
            I => prescaler_1_cry_3
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__7581\,
            I => \N__7577\
        );

    \I__1099\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7574\
        );

    \I__1098\ : InMux
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__7574\,
            I => \prescalerZ0Z_5\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__7571\,
            I => \prescalerZ0Z_5\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7566\,
            I => prescaler_1_cry_4
        );

    \I__1094\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7559\
        );

    \I__1093\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7556\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__7559\,
            I => \prescalerZ0Z_6\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__7556\,
            I => \prescalerZ0Z_6\
        );

    \I__1090\ : InMux
    port map (
            O => \N__7551\,
            I => prescaler_1_cry_5
        );

    \I__1089\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7544\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7541\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__7544\,
            I => \prescalerZ0Z_7\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__7541\,
            I => \prescalerZ0Z_7\
        );

    \I__1085\ : InMux
    port map (
            O => \N__7536\,
            I => prescaler_1_cry_6
        );

    \I__1084\ : InMux
    port map (
            O => \N__7533\,
            I => prescaler_1_cry_7
        );

    \I__1083\ : InMux
    port map (
            O => \N__7530\,
            I => \bfn_8_16_0_\
        );

    \I__1082\ : InMux
    port map (
            O => \N__7527\,
            I => \a.count_1_cry_20\
        );

    \I__1081\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7520\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7517\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__7520\,
            I => \N__7514\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__7517\,
            I => \a.countZ0Z_22\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__7514\,
            I => \a.countZ0Z_22\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7509\,
            I => \a.count_1_cry_21\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7502\
        );

    \I__1074\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7499\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__7502\,
            I => \a.countZ0Z_23\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__7499\,
            I => \a.countZ0Z_23\
        );

    \I__1071\ : InMux
    port map (
            O => \N__7494\,
            I => \a.count_1_cry_22\
        );

    \I__1070\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7487\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7484\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__7487\,
            I => \a.countZ0Z_24\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__7484\,
            I => \a.countZ0Z_24\
        );

    \I__1066\ : InMux
    port map (
            O => \N__7479\,
            I => \a.count_1_cry_23\
        );

    \I__1065\ : InMux
    port map (
            O => \N__7476\,
            I => \bfn_8_14_0_\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__7473\,
            I => \N__7469\
        );

    \I__1063\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__1062\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__7466\,
            I => \a.countZ0Z_25\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__7463\,
            I => \a.countZ0Z_25\
        );

    \I__1059\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7454\
        );

    \I__1058\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7451\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7454\,
            I => \a.countZ0Z_18\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__7451\,
            I => \a.countZ0Z_18\
        );

    \I__1055\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7442\
        );

    \I__1054\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7439\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7436\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__7439\,
            I => \a.countZ0Z_21\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__7436\,
            I => \a.countZ0Z_21\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__7431\,
            I => \N__7427\
        );

    \I__1049\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7424\
        );

    \I__1048\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7421\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__7424\,
            I => \a.countZ0Z_20\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__7421\,
            I => \a.countZ0Z_20\
        );

    \I__1045\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7412\
        );

    \I__1044\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7409\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__7412\,
            I => \a.countZ0Z_19\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__7409\,
            I => \a.countZ0Z_19\
        );

    \I__1041\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7401\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__7401\,
            I => \a.BUZZER3_15\
        );

    \I__1039\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7394\
        );

    \I__1038\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7391\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__7394\,
            I => \a.countZ0Z_12\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__7391\,
            I => \a.countZ0Z_12\
        );

    \I__1035\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7383\,
            I => \a.count_1_12\
        );

    \I__1033\ : InMux
    port map (
            O => \N__7380\,
            I => \a.count_1_cry_11\
        );

    \I__1032\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7373\
        );

    \I__1031\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7370\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__7373\,
            I => \a.countZ0Z_13\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__7370\,
            I => \a.countZ0Z_13\
        );

    \I__1028\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7362\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7362\,
            I => \a.count_1_13\
        );

    \I__1026\ : InMux
    port map (
            O => \N__7359\,
            I => \a.count_1_cry_12\
        );

    \I__1025\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7352\
        );

    \I__1024\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7349\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__7352\,
            I => \a.countZ0Z_14\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__7349\,
            I => \a.countZ0Z_14\
        );

    \I__1021\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__7341\,
            I => \a.count_1_14\
        );

    \I__1019\ : InMux
    port map (
            O => \N__7338\,
            I => \a.count_1_cry_13\
        );

    \I__1018\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7331\
        );

    \I__1017\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7328\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__7331\,
            I => \a.countZ0Z_15\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__7328\,
            I => \a.countZ0Z_15\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7323\,
            I => \a.count_1_cry_14\
        );

    \I__1013\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7316\
        );

    \I__1012\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7313\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__7316\,
            I => \a.countZ0Z_16\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__7313\,
            I => \a.countZ0Z_16\
        );

    \I__1009\ : InMux
    port map (
            O => \N__7308\,
            I => \a.count_1_cry_15\
        );

    \I__1008\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7301\
        );

    \I__1007\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7298\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__7301\,
            I => \a.countZ0Z_17\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__7298\,
            I => \a.countZ0Z_17\
        );

    \I__1004\ : InMux
    port map (
            O => \N__7293\,
            I => \bfn_8_13_0_\
        );

    \I__1003\ : InMux
    port map (
            O => \N__7290\,
            I => \a.count_1_cry_17\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7287\,
            I => \a.count_1_cry_18\
        );

    \I__1001\ : InMux
    port map (
            O => \N__7284\,
            I => \a.count_1_cry_19\
        );

    \I__1000\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7277\
        );

    \I__999\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7274\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__7277\,
            I => \a.countZ0Z_4\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__7274\,
            I => \a.countZ0Z_4\
        );

    \I__996\ : InMux
    port map (
            O => \N__7269\,
            I => \a.count_1_cry_3\
        );

    \I__995\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7262\
        );

    \I__994\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__7262\,
            I => \a.countZ0Z_5\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__7259\,
            I => \a.countZ0Z_5\
        );

    \I__991\ : InMux
    port map (
            O => \N__7254\,
            I => \a.count_1_cry_4\
        );

    \I__990\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7247\
        );

    \I__989\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7244\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__7247\,
            I => \a.countZ0Z_6\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__7244\,
            I => \a.countZ0Z_6\
        );

    \I__986\ : InMux
    port map (
            O => \N__7239\,
            I => \a.count_1_cry_5\
        );

    \I__985\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7232\
        );

    \I__984\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7229\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__7232\,
            I => \a.countZ0Z_7\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__7229\,
            I => \a.countZ0Z_7\
        );

    \I__981\ : InMux
    port map (
            O => \N__7224\,
            I => \a.count_1_cry_6\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__979\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__7215\,
            I => \N__7211\
        );

    \I__977\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7208\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__7211\,
            I => \a.countZ0Z_8\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__7208\,
            I => \a.countZ0Z_8\
        );

    \I__974\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__7200\,
            I => \a.count_1_8\
        );

    \I__972\ : InMux
    port map (
            O => \N__7197\,
            I => \a.count_1_cry_7\
        );

    \I__971\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7190\
        );

    \I__970\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7187\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__7190\,
            I => \a.countZ0Z_9\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__7187\,
            I => \a.countZ0Z_9\
        );

    \I__967\ : InMux
    port map (
            O => \N__7182\,
            I => \bfn_8_12_0_\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__7179\,
            I => \N__7176\
        );

    \I__965\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7172\
        );

    \I__964\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7169\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__7172\,
            I => \a.countZ0Z_10\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__7169\,
            I => \a.countZ0Z_10\
        );

    \I__961\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__7161\,
            I => \a.count_1_10\
        );

    \I__959\ : InMux
    port map (
            O => \N__7158\,
            I => \a.count_1_cry_9\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__957\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7148\
        );

    \I__956\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7145\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__7148\,
            I => \a.countZ0Z_11\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__7145\,
            I => \a.countZ0Z_11\
        );

    \I__953\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__7137\,
            I => \a.count_1_11\
        );

    \I__951\ : InMux
    port map (
            O => \N__7134\,
            I => \a.count_1_cry_10\
        );

    \I__950\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7127\
        );

    \I__949\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7124\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7121\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__7124\,
            I => \d1.countZ0Z_14\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__7121\,
            I => \d1.countZ0Z_14\
        );

    \I__945\ : InMux
    port map (
            O => \N__7116\,
            I => \d1.un3_count_cry_13\
        );

    \I__944\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7108\
        );

    \I__943\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7103\
        );

    \I__942\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7103\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__7108\,
            I => \d1.countZ0Z_15\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7103\,
            I => \d1.countZ0Z_15\
        );

    \I__939\ : InMux
    port map (
            O => \N__7098\,
            I => \d1.un3_count_cry_14\
        );

    \I__938\ : InMux
    port map (
            O => \N__7095\,
            I => \d1.un3_count_cry_15\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__7092\,
            I => \N__7087\
        );

    \I__936\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7084\
        );

    \I__935\ : InMux
    port map (
            O => \N__7090\,
            I => \N__7079\
        );

    \I__934\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7079\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7084\,
            I => \d1.countZ0Z_16\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7079\,
            I => \d1.countZ0Z_16\
        );

    \I__931\ : SRMux
    port map (
            O => \N__7074\,
            I => \N__7062\
        );

    \I__930\ : SRMux
    port map (
            O => \N__7073\,
            I => \N__7062\
        );

    \I__929\ : SRMux
    port map (
            O => \N__7072\,
            I => \N__7062\
        );

    \I__928\ : SRMux
    port map (
            O => \N__7071\,
            I => \N__7062\
        );

    \I__927\ : GlobalMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__926\ : gio2CtrlBuf
    port map (
            O => \N__7059\,
            I => \d1.idle_i_g\
        );

    \I__925\ : InMux
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__7047\,
            I => \N__7044\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__7044\,
            I => switch_dn_c
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__7041\,
            I => \N__7037\
        );

    \I__919\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7033\
        );

    \I__918\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7030\
        );

    \I__917\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7027\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__7033\,
            I => \a.countZ0Z_1\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7030\,
            I => \a.countZ0Z_1\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7027\,
            I => \a.countZ0Z_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7016\
        );

    \I__912\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7013\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__7016\,
            I => \a.countZ0Z_2\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__7013\,
            I => \a.countZ0Z_2\
        );

    \I__909\ : InMux
    port map (
            O => \N__7008\,
            I => \a.count_1_cry_1\
        );

    \I__908\ : InMux
    port map (
            O => \N__7005\,
            I => \N__7001\
        );

    \I__907\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6998\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__7001\,
            I => \a.countZ0Z_3\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6998\,
            I => \a.countZ0Z_3\
        );

    \I__904\ : InMux
    port map (
            O => \N__6993\,
            I => \a.count_1_cry_2\
        );

    \I__903\ : InMux
    port map (
            O => \N__6990\,
            I => \d1.un3_count_cry_4\
        );

    \I__902\ : InMux
    port map (
            O => \N__6987\,
            I => \d1.un3_count_cry_5\
        );

    \I__901\ : InMux
    port map (
            O => \N__6984\,
            I => \d1.un3_count_cry_6\
        );

    \I__900\ : InMux
    port map (
            O => \N__6981\,
            I => \d1.un3_count_cry_7\
        );

    \I__899\ : InMux
    port map (
            O => \N__6978\,
            I => \bfn_7_17_0_\
        );

    \I__898\ : InMux
    port map (
            O => \N__6975\,
            I => \d1.un3_count_cry_9\
        );

    \I__897\ : InMux
    port map (
            O => \N__6972\,
            I => \d1.un3_count_cry_10\
        );

    \I__896\ : InMux
    port map (
            O => \N__6969\,
            I => \d1.un3_count_cry_11\
        );

    \I__895\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6962\
        );

    \I__894\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__6959\,
            I => \d1.countZ0Z_13\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__6956\,
            I => \d1.countZ0Z_13\
        );

    \I__890\ : InMux
    port map (
            O => \N__6951\,
            I => \d1.un3_count_cry_12\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__888\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6941\
        );

    \I__887\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6938\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__6941\,
            I => \N__6935\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__6938\,
            I => \d1.syncZ0Z_1\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__6935\,
            I => \d1.syncZ0Z_1\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__6930\,
            I => \d1.trans_up_1_12_cascade_\
        );

    \I__882\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__6924\,
            I => \d1.g1_3\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__6921\,
            I => \d1.g1_4_cascade_\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__6918\,
            I => \N__6914\
        );

    \I__878\ : InMux
    port map (
            O => \N__6917\,
            I => \N__6909\
        );

    \I__877\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6906\
        );

    \I__876\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6901\
        );

    \I__875\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6901\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__6909\,
            I => \d1.countZ0Z_1\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__6906\,
            I => \d1.countZ0Z_1\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6901\,
            I => \d1.countZ0Z_1\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__6894\,
            I => \N__6890\
        );

    \I__870\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6886\
        );

    \I__869\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6881\
        );

    \I__868\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6881\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__6886\,
            I => \d1.countZ0Z_2\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__6881\,
            I => \d1.countZ0Z_2\
        );

    \I__865\ : InMux
    port map (
            O => \N__6876\,
            I => \d1.un3_count_cry_1\
        );

    \I__864\ : InMux
    port map (
            O => \N__6873\,
            I => \d1.un3_count_cry_2\
        );

    \I__863\ : InMux
    port map (
            O => \N__6870\,
            I => \d1.un3_count_cry_3\
        );

    \I__862\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6849\
        );

    \I__861\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6849\
        );

    \I__860\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6849\
        );

    \I__859\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6849\
        );

    \I__858\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6849\
        );

    \I__857\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6849\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6849\,
            I => \a.BUZZER3_20\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__6846\,
            I => \N__6837\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__6845\,
            I => \N__6834\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__6844\,
            I => \N__6831\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__6843\,
            I => \N__6828\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__6842\,
            I => \N__6825\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__6841\,
            I => \N__6822\
        );

    \I__849\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6819\
        );

    \I__848\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6810\
        );

    \I__847\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6810\
        );

    \I__846\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6810\
        );

    \I__845\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6810\
        );

    \I__844\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6805\
        );

    \I__843\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6805\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__6819\,
            I => \a.BUZZER3_19\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__6810\,
            I => \a.BUZZER3_19\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6805\,
            I => \a.BUZZER3_19\
        );

    \I__839\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6795\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__6795\,
            I => \a.BUZZER3_18\
        );

    \I__837\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6789\,
            I => \a.BUZZER3_17\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__6786\,
            I => \a.BUZZER3_16_cascade_\
        );

    \I__834\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__6780\,
            I => \N__6771\
        );

    \I__832\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6758\
        );

    \I__831\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6758\
        );

    \I__830\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6758\
        );

    \I__829\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6758\
        );

    \I__828\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6758\
        );

    \I__827\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6758\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__6771\,
            I => \a.BUZZER3_24\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__6758\,
            I => \a.BUZZER3_24\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__6753\,
            I => \a.BUZZER3_14_cascade_\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__6750\,
            I => \a.BUZZER3_20_cascade_\
        );

    \I__822\ : IoInMux
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__820\ : Span12Mux_s10_h
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__819\ : Span12Mux_v
    port map (
            O => \N__6738\,
            I => \N__6734\
        );

    \I__818\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6731\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__6734\,
            I => \BUZZER_c\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__6731\,
            I => \BUZZER_c\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__814\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6719\
        );

    \I__813\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6716\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6713\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__6716\,
            I => \display1.prescalerZ0Z_22\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__6713\,
            I => \display1.prescalerZ0Z_22\
        );

    \I__809\ : InMux
    port map (
            O => \N__6708\,
            I => \display1.prescaler_2_cry_21\
        );

    \I__808\ : InMux
    port map (
            O => \N__6705\,
            I => \display1.prescaler_2_cry_22\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__806\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6696\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6696\,
            I => \N__6692\
        );

    \I__804\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6689\
        );

    \I__803\ : Span4Mux_h
    port map (
            O => \N__6692\,
            I => \N__6686\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__6689\,
            I => \display1.prescalerZ0Z_23\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__6686\,
            I => \display1.prescalerZ0Z_23\
        );

    \I__800\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6677\
        );

    \I__799\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6674\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6677\,
            I => \display1.prescalerZ0Z_12\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__6674\,
            I => \display1.prescalerZ0Z_12\
        );

    \I__796\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6665\
        );

    \I__795\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6662\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6665\,
            I => \display1.prescalerZ0Z_11\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__6662\,
            I => \display1.prescalerZ0Z_11\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__6657\,
            I => \N__6653\
        );

    \I__791\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6650\
        );

    \I__790\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6647\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6650\,
            I => \display1.prescalerZ0Z_13\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__6647\,
            I => \display1.prescalerZ0Z_13\
        );

    \I__787\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6638\
        );

    \I__786\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6635\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__6638\,
            I => \display1.prescalerZ0Z_10\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__6635\,
            I => \display1.prescalerZ0Z_10\
        );

    \I__783\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__6621\,
            I => \display1.prescaler8_12\
        );

    \I__779\ : IoInMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__777\ : Span12Mux_s9_h
    port map (
            O => \N__6612\,
            I => \N__6609\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__6609\,
            I => \d1.idle_i\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__6606\,
            I => \d1.trans_up_1_11_cascade_\
        );

    \I__774\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6596\
        );

    \I__772\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6593\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__6596\,
            I => \display1.prescalerZ0Z_14\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__6593\,
            I => \display1.prescalerZ0Z_14\
        );

    \I__769\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6585\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__6582\,
            I => \display1.prescaler_2_14\
        );

    \I__766\ : InMux
    port map (
            O => \N__6579\,
            I => \display1.prescaler_2_cry_13\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__6576\,
            I => \N__6572\
        );

    \I__764\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6569\
        );

    \I__763\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6566\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__6569\,
            I => \N__6563\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__6566\,
            I => \N__6560\
        );

    \I__760\ : Odrv12
    port map (
            O => \N__6563\,
            I => \display1.prescalerZ0Z_15\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__6560\,
            I => \display1.prescalerZ0Z_15\
        );

    \I__758\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__6552\,
            I => \N__6549\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__6549\,
            I => \display1.prescaler_2_15\
        );

    \I__755\ : InMux
    port map (
            O => \N__6546\,
            I => \display1.prescaler_2_cry_14\
        );

    \I__754\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6539\
        );

    \I__753\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6536\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6533\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__6536\,
            I => \display1.prescalerZ0Z_16\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__6533\,
            I => \display1.prescalerZ0Z_16\
        );

    \I__749\ : InMux
    port map (
            O => \N__6528\,
            I => \display1.prescaler_2_cry_15\
        );

    \I__748\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6521\
        );

    \I__747\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6518\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__6518\,
            I => \N__6510\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__6515\,
            I => \N__6510\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__6510\,
            I => \display1.prescalerZ0Z_17\
        );

    \I__742\ : InMux
    port map (
            O => \N__6507\,
            I => \bfn_5_15_0_\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__740\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__6498\,
            I => \N__6494\
        );

    \I__738\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6491\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__6494\,
            I => \N__6488\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__6491\,
            I => \display1.prescalerZ0Z_18\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__6488\,
            I => \display1.prescalerZ0Z_18\
        );

    \I__734\ : InMux
    port map (
            O => \N__6483\,
            I => \display1.prescaler_2_cry_17\
        );

    \I__733\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6476\
        );

    \I__732\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6473\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6470\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__6473\,
            I => \display1.prescalerZ0Z_19\
        );

    \I__729\ : Odrv4
    port map (
            O => \N__6470\,
            I => \display1.prescalerZ0Z_19\
        );

    \I__728\ : InMux
    port map (
            O => \N__6465\,
            I => \display1.prescaler_2_cry_18\
        );

    \I__727\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6458\
        );

    \I__726\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6455\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__6458\,
            I => \N__6452\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__6455\,
            I => \display1.prescalerZ0Z_20\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__6452\,
            I => \display1.prescalerZ0Z_20\
        );

    \I__722\ : InMux
    port map (
            O => \N__6447\,
            I => \display1.prescaler_2_cry_19\
        );

    \I__721\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6440\
        );

    \I__720\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6437\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__6440\,
            I => \N__6434\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__6437\,
            I => \display1.prescalerZ0Z_21\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__6434\,
            I => \display1.prescalerZ0Z_21\
        );

    \I__716\ : InMux
    port map (
            O => \N__6429\,
            I => \display1.prescaler_2_cry_20\
        );

    \I__715\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6419\
        );

    \I__713\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6416\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__6419\,
            I => \display1.prescalerZ0Z_6\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__6416\,
            I => \display1.prescalerZ0Z_6\
        );

    \I__710\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__6405\,
            I => \display1.prescaler_2_6\
        );

    \I__707\ : InMux
    port map (
            O => \N__6402\,
            I => \display1.prescaler_2_cry_5\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__6399\,
            I => \N__6395\
        );

    \I__705\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6392\
        );

    \I__704\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6389\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__6392\,
            I => \display1.prescalerZ0Z_7\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__6389\,
            I => \display1.prescalerZ0Z_7\
        );

    \I__701\ : InMux
    port map (
            O => \N__6384\,
            I => \display1.prescaler_2_cry_6\
        );

    \I__700\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6374\
        );

    \I__698\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6371\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__6374\,
            I => \display1.prescalerZ0Z_8\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__6371\,
            I => \display1.prescalerZ0Z_8\
        );

    \I__695\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6363\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__6360\,
            I => \display1.prescaler_2_8\
        );

    \I__692\ : InMux
    port map (
            O => \N__6357\,
            I => \display1.prescaler_2_cry_7\
        );

    \I__691\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__6351\,
            I => \N__6347\
        );

    \I__689\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6344\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__6347\,
            I => \display1.prescalerZ0Z_9\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__6344\,
            I => \display1.prescalerZ0Z_9\
        );

    \I__686\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6336\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__6333\,
            I => \display1.prescaler_2_9\
        );

    \I__683\ : InMux
    port map (
            O => \N__6330\,
            I => \bfn_5_14_0_\
        );

    \I__682\ : InMux
    port map (
            O => \N__6327\,
            I => \display1.prescaler_2_cry_9\
        );

    \I__681\ : InMux
    port map (
            O => \N__6324\,
            I => \display1.prescaler_2_cry_10\
        );

    \I__680\ : InMux
    port map (
            O => \N__6321\,
            I => \display1.prescaler_2_cry_11\
        );

    \I__679\ : InMux
    port map (
            O => \N__6318\,
            I => \display1.prescaler_2_cry_12\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__6315\,
            I => \display1.prescaler8_17_cascade_\
        );

    \I__677\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6298\
        );

    \I__676\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6298\
        );

    \I__675\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6298\
        );

    \I__674\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6291\
        );

    \I__673\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6291\
        );

    \I__672\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6291\
        );

    \I__671\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6286\
        );

    \I__670\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6286\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__6298\,
            I => \display1.prescaler8_21\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__6291\,
            I => \display1.prescaler8_21\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__6286\,
            I => \display1.prescaler8_21\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__6279\,
            I => \N__6274\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__6278\,
            I => \N__6268\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__6277\,
            I => \N__6265\
        );

    \I__663\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6256\
        );

    \I__662\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6256\
        );

    \I__661\ : InMux
    port map (
            O => \N__6272\,
            I => \N__6256\
        );

    \I__660\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6256\
        );

    \I__659\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6249\
        );

    \I__658\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6249\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6246\
        );

    \I__656\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6241\
        );

    \I__655\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6241\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__6249\,
            I => \display1.prescaler8_17\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__6246\,
            I => \display1.prescaler8_17\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__6241\,
            I => \display1.prescaler8_17\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__6234\,
            I => \N__6230\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__6233\,
            I => \N__6227\
        );

    \I__649\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6215\
        );

    \I__648\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6215\
        );

    \I__647\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6215\
        );

    \I__646\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6212\
        );

    \I__645\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6205\
        );

    \I__644\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6205\
        );

    \I__643\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6205\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6198\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__6212\,
            I => \N__6198\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6195\
        );

    \I__639\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6190\
        );

    \I__638\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6190\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__6198\,
            I => \display1.prescaler8_16\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__6195\,
            I => \display1.prescaler8_16\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__6190\,
            I => \display1.prescaler8_16\
        );

    \I__634\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6180\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6180\,
            I => \N__6177\
        );

    \I__632\ : Span4Mux_h
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__6174\,
            I => \display1.prescaler8_13\
        );

    \I__630\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6163\
        );

    \I__628\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6158\
        );

    \I__627\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6158\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__6163\,
            I => \display1.prescalerZ0Z_1\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__6158\,
            I => \display1.prescalerZ0Z_1\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__623\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6144\
        );

    \I__622\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6139\
        );

    \I__621\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6139\
        );

    \I__620\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6136\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6133\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__6139\,
            I => \display1.prescalerZ0Z_0\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__6136\,
            I => \display1.prescalerZ0Z_0\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__6133\,
            I => \display1.prescalerZ0Z_0\
        );

    \I__615\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6122\
        );

    \I__614\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6119\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__6122\,
            I => \display1.prescalerZ0Z_2\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__6119\,
            I => \display1.prescalerZ0Z_2\
        );

    \I__611\ : InMux
    port map (
            O => \N__6114\,
            I => \display1.prescaler_2_cry_1\
        );

    \I__610\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6107\
        );

    \I__609\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6104\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__6107\,
            I => \display1.prescalerZ0Z_3\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__6104\,
            I => \display1.prescalerZ0Z_3\
        );

    \I__606\ : InMux
    port map (
            O => \N__6099\,
            I => \display1.prescaler_2_cry_2\
        );

    \I__605\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6093\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__6093\,
            I => \N__6089\
        );

    \I__603\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6086\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__6089\,
            I => \display1.prescalerZ0Z_4\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__6086\,
            I => \display1.prescalerZ0Z_4\
        );

    \I__600\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__6078\,
            I => \N__6075\
        );

    \I__598\ : Span4Mux_h
    port map (
            O => \N__6075\,
            I => \N__6072\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__6072\,
            I => \display1.prescaler_2_4\
        );

    \I__596\ : InMux
    port map (
            O => \N__6069\,
            I => \display1.prescaler_2_cry_3\
        );

    \I__595\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6062\
        );

    \I__594\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6059\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__6062\,
            I => \display1.prescalerZ0Z_5\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__6059\,
            I => \display1.prescalerZ0Z_5\
        );

    \I__591\ : InMux
    port map (
            O => \N__6054\,
            I => \display1.prescaler_2_cry_4\
        );

    \I__590\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__6048\,
            I => \display1.prescaler8_14\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__6045\,
            I => \display1.prescaler8_15_cascade_\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__6042\,
            I => \display1.prescaler8_21_cascade_\
        );

    \I__586\ : IoInMux
    port map (
            O => \N__6039\,
            I => \N__6036\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__6036\,
            I => \N__6033\
        );

    \I__584\ : Span12Mux_s4_h
    port map (
            O => \N__6033\,
            I => \N__6030\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__6030\,
            I => \SEG1_c_2\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__6027\,
            I => \N__6024\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__6024\,
            I => \N__6021\
        );

    \I__580\ : IoSpan4Mux
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__579\ : Span4Mux_s3_v
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__6009\,
            I => \SEG1_c_0\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__6006\,
            I => \display1.prescaler8_cascade_\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__6003\,
            I => \N__5997\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__6002\,
            I => \N__5994\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__6001\,
            I => \N__5990\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__6000\,
            I => \N__5987\
        );

    \I__570\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5977\
        );

    \I__569\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5977\
        );

    \I__568\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5977\
        );

    \I__567\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5968\
        );

    \I__566\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5968\
        );

    \I__565\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5968\
        );

    \I__564\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5968\
        );

    \I__563\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5965\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5977\,
            I => \display1.digit_dataZ0Z_3\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5968\,
            I => \display1.digit_dataZ0Z_3\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5965\,
            I => \display1.digit_dataZ0Z_3\
        );

    \I__559\ : IoInMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__557\ : IoSpan4Mux
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__556\ : Span4Mux_s3_h
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__5940\,
            I => \DIGIT_c_0\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__5937\,
            I => \N__5932\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__5936\,
            I => \N__5927\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__5935\,
            I => \N__5922\
        );

    \I__549\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5913\
        );

    \I__548\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5913\
        );

    \I__547\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5913\
        );

    \I__546\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5913\
        );

    \I__545\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5906\
        );

    \I__544\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5906\
        );

    \I__543\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5906\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5913\,
            I => \display1.digit_dataZ0Z_2\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__5906\,
            I => \display1.digit_dataZ0Z_2\
        );

    \I__540\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5886\
        );

    \I__539\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5886\
        );

    \I__538\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5886\
        );

    \I__537\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5886\
        );

    \I__536\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5879\
        );

    \I__535\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5879\
        );

    \I__534\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5879\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5886\,
            I => \display1.digit_dataZ0Z_1\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5879\,
            I => \display1.digit_dataZ0Z_1\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__5874\,
            I => \N__5866\
        );

    \I__530\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5863\
        );

    \I__529\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5854\
        );

    \I__528\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5854\
        );

    \I__527\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5854\
        );

    \I__526\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5854\
        );

    \I__525\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5851\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__5863\,
            I => \display1.digit_posnZ0\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5854\,
            I => \display1.digit_posnZ0\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__5851\,
            I => \display1.digit_posnZ0\
        );

    \I__521\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5829\
        );

    \I__520\ : InMux
    port map (
            O => \N__5843\,
            I => \N__5829\
        );

    \I__519\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5829\
        );

    \I__518\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5829\
        );

    \I__517\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5822\
        );

    \I__516\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5822\
        );

    \I__515\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5822\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5829\,
            I => \display1.digit_dataZ0Z_0\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__5822\,
            I => \display1.digit_dataZ0Z_0\
        );

    \I__512\ : CEMux
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5814\,
            I => \display1.prescaler8\
        );

    \I__510\ : IoInMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__508\ : IoSpan4Mux
    port map (
            O => \N__5805\,
            I => \N__5802\
        );

    \I__507\ : Span4Mux_s1_h
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__5799\,
            I => \SEG1_c_5\
        );

    \I__505\ : IoInMux
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__5793\,
            I => \N__5790\
        );

    \I__503\ : IoSpan4Mux
    port map (
            O => \N__5790\,
            I => \N__5787\
        );

    \I__502\ : Span4Mux_s3_h
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__5784\,
            I => \SEG1_c_6\
        );

    \I__500\ : IoInMux
    port map (
            O => \N__5781\,
            I => \N__5778\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__5775\,
            I => \SEG1_c_4\
        );

    \I__497\ : IoInMux
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5766\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__5766\,
            I => \SEG1_c_3\
        );

    \I__494\ : IoInMux
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__492\ : Span4Mux_s3_h
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__5754\,
            I => \N__5751\
        );

    \I__490\ : Odrv4
    port map (
            O => \N__5751\,
            I => \SEG1_c_1\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => prescaler_1_cry_8,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => prescaler_1_cry_16,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => prescaler_1_cry_24,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \display2.prescaler_2_cry_8\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \display2.prescaler_2_cry_16\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \display1.prescaler_2_cry_8\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \display1.prescaler_2_cry_16\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d4.un3_count_cry_8\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d3.un3_count_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d2.un3_count_cry_8\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d1.un3_count_cry_8\,
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \a.count_1_cry_8\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \a.count_1_cry_16\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \a.count_1_cry_24\,
            carryinitout => \bfn_8_14_0_\
        );

    \un1_state_3_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10560\,
            GLOBALBUFFEROUTPUT => un1_state_3_g
        );

    \d4.sync_1_RNIQPEK_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8529\,
            GLOBALBUFFEROUTPUT => \d4.idle_i_g\
        );

    \d3.state_RNIOCAC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12543\,
            GLOBALBUFFEROUTPUT => \d3.idle_i_g\
        );

    \d2.sync_1_RNIMV5K_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11928\,
            GLOBALBUFFEROUTPUT => \d2.idle_i_g\
        );

    \d1.sync_1_RNIKI1C_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6618\,
            GLOBALBUFFEROUTPUT => \d1.idle_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \display1.decoder.SEG_5_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100111111"
        )
    port map (
            in0 => \N__5843\,
            in1 => \N__5900\,
            in2 => \N__6001\,
            in3 => \N__5931\,
            lcout => \SEG1_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_6_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011000100111"
        )
    port map (
            in0 => \N__5901\,
            in1 => \N__5986\,
            in2 => \N__5937\,
            in3 => \N__5844\,
            lcout => \SEG1_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_4_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100111011"
        )
    port map (
            in0 => \N__5842\,
            in1 => \N__5899\,
            in2 => \N__6000\,
            in3 => \N__5930\,
            lcout => \SEG1_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_3_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000100111"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__5985\,
            in2 => \N__5936\,
            in3 => \N__5841\,
            lcout => \SEG1_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_1_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100110001"
        )
    port map (
            in0 => \N__5839\,
            in1 => \N__5896\,
            in2 => \N__6002\,
            in3 => \N__5925\,
            lcout => \SEG1_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_2_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000010101"
        )
    port map (
            in0 => \N__5840\,
            in1 => \N__5897\,
            in2 => \N__6003\,
            in3 => \N__5926\,
            lcout => \SEG1_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.decoder.SEG_0_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000110110"
        )
    port map (
            in0 => \N__5895\,
            in1 => \N__5993\,
            in2 => \N__5935\,
            in3 => \N__5838\,
            lcout => \SEG1_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNI2HUD5_16_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__6203\,
            in2 => \_gnd_net_\,
            in3 => \N__6305\,
            lcout => \display1.prescaler8\,
            ltout => \display1.prescaler8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.digit_data_3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__5873\,
            in1 => \N__5984\,
            in2 => \N__6006\,
            in3 => \N__10407\,
            lcout => \display1.digit_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.digit_posn_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__6204\,
            in2 => \N__5874\,
            in3 => \N__6306\,
            lcout => \display1.digit_posnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.DIGIT_e_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5872\,
            lcout => \DIGIT_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14265\,
            ce => \N__5817\,
            sr => \_gnd_net_\
        );

    \display1.digit_data_e_0_2_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5871\,
            in1 => \N__10482\,
            in2 => \_gnd_net_\,
            in3 => \N__10600\,
            lcout => \display1.digit_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14265\,
            ce => \N__5817\,
            sr => \_gnd_net_\
        );

    \display1.digit_data_e_0_1_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10446\,
            in1 => \N__12507\,
            in2 => \_gnd_net_\,
            in3 => \N__5870\,
            lcout => \display1.digit_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14265\,
            ce => \N__5817\,
            sr => \_gnd_net_\
        );

    \display1.digit_data_e_0_0_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5869\,
            in1 => \N__10368\,
            in2 => \_gnd_net_\,
            in3 => \N__12456\,
            lcout => \display1.digit_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14265\,
            ce => \N__5817\,
            sr => \_gnd_net_\
        );

    \display1.prescaler_8_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6309\,
            in1 => \N__6273\,
            in2 => \N__6234\,
            in3 => \N__6366\,
            lcout => \display1.prescalerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_4_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6225\,
            in1 => \N__6081\,
            in2 => \N__6279\,
            in3 => \N__6307\,
            lcout => \display1.prescalerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNID8UQ_1_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6599\,
            in1 => \N__6350\,
            in2 => \N__6576\,
            in3 => \N__6166\,
            lcout => \display1.prescaler8_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNIVNSK_23_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6377\,
            in1 => \N__6422\,
            in2 => \N__6702\,
            in3 => \N__6092\,
            lcout => OPEN,
            ltout => \display1.prescaler8_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNIN1N53_1_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__6183\,
            in2 => \N__6045\,
            in3 => \N__6630\,
            lcout => \display1.prescaler8_21\,
            ltout => \display1.prescaler8_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_0_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__6271\,
            in1 => \N__6226\,
            in2 => \N__6042\,
            in3 => \N__6148\,
            lcout => \display1.prescalerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_6_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6308\,
            in1 => \N__6272\,
            in2 => \N__6233\,
            in3 => \N__6411\,
            lcout => \display1.prescalerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_1_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6149\,
            lcout => \display1.prescalerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_9_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6312\,
            in1 => \N__6224\,
            in2 => \N__6278\,
            in3 => \N__6339\,
            lcout => \display1.prescalerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNI0V011_16_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6525\,
            in1 => \N__6543\,
            in2 => \N__6504\,
            in3 => \N__6147\,
            lcout => \display1.prescaler8_17\,
            ltout => \display1.prescaler8_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_14_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6222\,
            in1 => \N__6588\,
            in2 => \N__6315\,
            in3 => \N__6310\,
            lcout => \display1.prescalerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_15_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__6223\,
            in2 => \N__6277\,
            in3 => \N__6555\,
            lcout => \display1.prescalerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNIBG671_19_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6444\,
            in1 => \N__6462\,
            in2 => \N__6726\,
            in3 => \N__6480\,
            lcout => \display1.prescaler8_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNI9TOE_2_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6065\,
            in1 => \N__6125\,
            in2 => \N__6399\,
            in3 => \N__6110\,
            lcout => \display1.prescaler8_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_2_cry_1_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6171\,
            in2 => \N__6153\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \display1.prescaler_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_2_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6126\,
            in2 => \_gnd_net_\,
            in3 => \N__6114\,
            lcout => \display1.prescalerZ0Z_2\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_1\,
            carryout => \display1.prescaler_2_cry_2\,
            clk => \N__14264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6111\,
            in2 => \_gnd_net_\,
            in3 => \N__6099\,
            lcout => \display1.prescalerZ0Z_3\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_2\,
            carryout => \display1.prescaler_2_cry_3\,
            clk => \N__14264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_4_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6096\,
            in2 => \_gnd_net_\,
            in3 => \N__6069\,
            lcout => \display1.prescaler_2_4\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_3\,
            carryout => \display1.prescaler_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_5_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6066\,
            in2 => \_gnd_net_\,
            in3 => \N__6054\,
            lcout => \display1.prescalerZ0Z_5\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_4\,
            carryout => \display1.prescaler_2_cry_5\,
            clk => \N__14264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6426\,
            in2 => \_gnd_net_\,
            in3 => \N__6402\,
            lcout => \display1.prescaler_2_6\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_5\,
            carryout => \display1.prescaler_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_7_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6398\,
            in2 => \_gnd_net_\,
            in3 => \N__6384\,
            lcout => \display1.prescalerZ0Z_7\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_6\,
            carryout => \display1.prescaler_2_cry_7\,
            clk => \N__14264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_8_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6381\,
            in2 => \_gnd_net_\,
            in3 => \N__6357\,
            lcout => \display1.prescaler_2_8\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_7\,
            carryout => \display1.prescaler_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_9_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6354\,
            in2 => \_gnd_net_\,
            in3 => \N__6330\,
            lcout => \display1.prescaler_2_9\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \display1.prescaler_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_10_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6642\,
            in2 => \_gnd_net_\,
            in3 => \N__6327\,
            lcout => \display1.prescalerZ0Z_10\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_9\,
            carryout => \display1.prescaler_2_cry_10\,
            clk => \N__14261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6669\,
            in2 => \_gnd_net_\,
            in3 => \N__6324\,
            lcout => \display1.prescalerZ0Z_11\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_10\,
            carryout => \display1.prescaler_2_cry_11\,
            clk => \N__14261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_12_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6681\,
            in2 => \_gnd_net_\,
            in3 => \N__6321\,
            lcout => \display1.prescalerZ0Z_12\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_11\,
            carryout => \display1.prescaler_2_cry_12\,
            clk => \N__14261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_13_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6656\,
            in2 => \_gnd_net_\,
            in3 => \N__6318\,
            lcout => \display1.prescalerZ0Z_13\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_12\,
            carryout => \display1.prescaler_2_cry_13\,
            clk => \N__14261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_14_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6603\,
            in2 => \_gnd_net_\,
            in3 => \N__6579\,
            lcout => \display1.prescaler_2_14\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_13\,
            carryout => \display1.prescaler_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNO_0_15_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6575\,
            in2 => \_gnd_net_\,
            in3 => \N__6546\,
            lcout => \display1.prescaler_2_15\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_14\,
            carryout => \display1.prescaler_2_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_16_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6542\,
            in2 => \_gnd_net_\,
            in3 => \N__6528\,
            lcout => \display1.prescalerZ0Z_16\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_15\,
            carryout => \display1.prescaler_2_cry_16\,
            clk => \N__14261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_17_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6524\,
            in2 => \_gnd_net_\,
            in3 => \N__6507\,
            lcout => \display1.prescalerZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \display1.prescaler_2_cry_17\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_18_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6497\,
            in2 => \_gnd_net_\,
            in3 => \N__6483\,
            lcout => \display1.prescalerZ0Z_18\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_17\,
            carryout => \display1.prescaler_2_cry_18\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_19_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6479\,
            in2 => \_gnd_net_\,
            in3 => \N__6465\,
            lcout => \display1.prescalerZ0Z_19\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_18\,
            carryout => \display1.prescaler_2_cry_19\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_20_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6461\,
            in2 => \_gnd_net_\,
            in3 => \N__6447\,
            lcout => \display1.prescalerZ0Z_20\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_19\,
            carryout => \display1.prescaler_2_cry_20\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_21_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6443\,
            in2 => \_gnd_net_\,
            in3 => \N__6429\,
            lcout => \display1.prescalerZ0Z_21\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_20\,
            carryout => \display1.prescaler_2_cry_21\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_22_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6722\,
            in2 => \_gnd_net_\,
            in3 => \N__6708\,
            lcout => \display1.prescalerZ0Z_22\,
            ltout => OPEN,
            carryin => \display1.prescaler_2_cry_21\,
            carryout => \display1.prescaler_2_cry_22\,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_23_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6695\,
            in2 => \_gnd_net_\,
            in3 => \N__6705\,
            lcout => \display1.prescalerZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display1.prescaler_RNI24371_10_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__6668\,
            in2 => \N__6657\,
            in3 => \N__6641\,
            lcout => \display1.prescaler8_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_RNIKI1C_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6944\,
            in2 => \_gnd_net_\,
            in3 => \N__9065\,
            lcout => \d1.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_stored_e_0_3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13899\,
            lcout => \mins_storedZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14252\,
            ce => \N__10774\,
            sr => \_gnd_net_\
        );

    \d1.count_1_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6917\,
            in2 => \_gnd_net_\,
            in3 => \N__8309\,
            lcout => \d1.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14245\,
            ce => 'H',
            sr => \N__7071\
        );

    \d1.count_RNI0AFK_0_16_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6913\,
            in1 => \N__7090\,
            in2 => \N__6894\,
            in3 => \N__7112\,
            lcout => \d1.g0_1_a5_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI0AFK_16_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7111\,
            in1 => \N__6889\,
            in2 => \N__7092\,
            in3 => \N__6912\,
            lcout => \d1.trans_up_1_11\,
            ltout => \d1.trans_up_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIRPKB1_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__9048\,
            in1 => \N__12798\,
            in2 => \N__6606\,
            in3 => \N__11902\,
            lcout => \d1.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.stateZ0_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9052\,
            in2 => \_gnd_net_\,
            in3 => \N__10221\,
            lcout => \d1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNIQ0UE1_22_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7005\,
            in1 => \N__7020\,
            in2 => \N__7041\,
            in3 => \N__7524\,
            lcout => OPEN,
            ltout => \a.BUZZER3_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNI7VOF2_4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10689\,
            in1 => \N__7281\,
            in2 => \N__6753\,
            in3 => \N__8662\,
            lcout => \a.BUZZER3_20\,
            ltout => \a.BUZZER3_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.BUZZER_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__6737\,
            in1 => \N__6840\,
            in2 => \N__6750\,
            in3 => \N__6783\,
            lcout => \BUZZER_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNI39TE1_10_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7236\,
            in1 => \N__7251\,
            in2 => \N__7179\,
            in3 => \N__7266\,
            lcout => \a.BUZZER3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_11_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6775\,
            in1 => \N__6863\,
            in2 => \N__6843\,
            in3 => \N__7140\,
            lcout => \a.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_10_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6862\,
            in1 => \N__6774\,
            in2 => \N__6841\,
            in3 => \N__7164\,
            lcout => \a.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_14_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6778\,
            in1 => \N__6866\,
            in2 => \N__6845\,
            in3 => \N__7344\,
            lcout => \a.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNIE4K61_11_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7376\,
            in1 => \N__7397\,
            in2 => \N__7155\,
            in3 => \N__7355\,
            lcout => \a.BUZZER3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_13_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6777\,
            in1 => \N__6865\,
            in2 => \N__6844\,
            in3 => \N__7365\,
            lcout => \a.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_8_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6779\,
            in1 => \N__6867\,
            in2 => \N__6846\,
            in3 => \N__7203\,
            lcout => \a.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_12_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6864\,
            in1 => \N__6776\,
            in2 => \N__6842\,
            in3 => \N__7386\,
            lcout => \a.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNIS97C1_23_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7505\,
            in1 => \N__7194\,
            in2 => \N__7221\,
            in3 => \N__7490\,
            lcout => \a.BUZZER3_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13917\,
            lcout => \d1.syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNISJL61_25_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7334\,
            in1 => \N__7304\,
            in2 => \N__7473\,
            in3 => \N__7319\,
            lcout => OPEN,
            ltout => \a.BUZZER3_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNIUI705_11_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6798\,
            in1 => \N__6792\,
            in2 => \N__6786\,
            in3 => \N__7404\,
            lcout => \a.BUZZER3_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7652\,
            lcout => \prescalerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14246\,
            ce => \N__8053\,
            sr => \_gnd_net_\
        );

    \prescaler_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7675\,
            lcout => \prescalerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14246\,
            ce => \N__8053\,
            sr => \_gnd_net_\
        );

    \d1.count_RNI2PCE_0_3_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11025\,
            in1 => \N__11052\,
            in2 => \N__11001\,
            in3 => \N__10968\,
            lcout => \d1.g0_1_a5_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI5QJP_11_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8611\,
            in1 => \N__8270\,
            in2 => \N__9066\,
            in3 => \N__8303\,
            lcout => \d1.g0_1_a5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_0_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8304\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \d1.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14238\,
            ce => 'H',
            sr => \N__7072\
        );

    \d1.count_RNI2PCE_3_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11026\,
            in1 => \N__11053\,
            in2 => \N__11002\,
            in3 => \N__10969\,
            lcout => \d1.trans_up_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_RNI5IAP_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__7131\,
            in1 => \N__9056\,
            in2 => \N__6948\,
            in3 => \N__6966\,
            lcout => \d1.trans_up_1_12\,
            ltout => \d1.trans_up_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI9D0D1_3_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__9167\,
            in1 => \_gnd_net_\,
            in2 => \N__6930\,
            in3 => \N__8331\,
            lcout => OPEN,
            ltout => \d1.g1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIINS67_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__6927\,
            in1 => \N__10167\,
            in2 => \N__6921\,
            in3 => \N__9126\,
            lcout => \d1.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.un3_count_cry_1_c_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8308\,
            in2 => \N__6918\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \d1.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6893\,
            in2 => \_gnd_net_\,
            in3 => \N__6876\,
            lcout => \d1.countZ0Z_2\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_1\,
            carryout => \d1.un3_count_cry_2\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_3_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10973\,
            in2 => \_gnd_net_\,
            in3 => \N__6873\,
            lcout => \d1.countZ0Z_3\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_2\,
            carryout => \d1.un3_count_cry_3\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_4_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11030\,
            in2 => \_gnd_net_\,
            in3 => \N__6870\,
            lcout => \d1.countZ0Z_4\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_3\,
            carryout => \d1.un3_count_cry_4\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_5_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11057\,
            in2 => \_gnd_net_\,
            in3 => \N__6990\,
            lcout => \d1.countZ0Z_5\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_4\,
            carryout => \d1.un3_count_cry_5\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_6_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11006\,
            in2 => \_gnd_net_\,
            in3 => \N__6987\,
            lcout => \d1.countZ0Z_6\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_5\,
            carryout => \d1.un3_count_cry_6\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_7_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8876\,
            in2 => \_gnd_net_\,
            in3 => \N__6984\,
            lcout => \d1.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_6\,
            carryout => \d1.un3_count_cry_7\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_8_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8929\,
            in2 => \_gnd_net_\,
            in3 => \N__6981\,
            lcout => \d1.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_7\,
            carryout => \d1.un3_count_cry_8\,
            clk => \N__14232\,
            ce => 'H',
            sr => \N__7073\
        );

    \d1.count_9_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8956\,
            in2 => \_gnd_net_\,
            in3 => \N__6978\,
            lcout => \d1.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \d1.un3_count_cry_9\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_10_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8899\,
            in2 => \_gnd_net_\,
            in3 => \N__6975\,
            lcout => \d1.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_9\,
            carryout => \d1.un3_count_cry_10\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_11_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8269\,
            in2 => \_gnd_net_\,
            in3 => \N__6972\,
            lcout => \d1.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_10\,
            carryout => \d1.un3_count_cry_11\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_12_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8610\,
            in2 => \_gnd_net_\,
            in3 => \N__6969\,
            lcout => \d1.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_11\,
            carryout => \d1.un3_count_cry_12\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_13_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6965\,
            in2 => \_gnd_net_\,
            in3 => \N__6951\,
            lcout => \d1.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_12\,
            carryout => \d1.un3_count_cry_13\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_14_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7130\,
            in2 => \_gnd_net_\,
            in3 => \N__7116\,
            lcout => \d1.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_13\,
            carryout => \d1.un3_count_cry_14\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_15_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7113\,
            in2 => \_gnd_net_\,
            in3 => \N__7098\,
            lcout => \d1.countZ0Z_15\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_14\,
            carryout => \d1.un3_count_cry_15\,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d1.count_16_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7091\,
            in2 => \_gnd_net_\,
            in3 => \N__7095\,
            lcout => \d1.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14224\,
            ce => 'H',
            sr => \N__7074\
        );

    \d2.sync_0_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \d2.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8664\,
            in2 => \_gnd_net_\,
            in3 => \N__7040\,
            lcout => \a.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_1_cry_1_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7036\,
            in2 => \N__8663\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \a.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7019\,
            in2 => \_gnd_net_\,
            in3 => \N__7008\,
            lcout => \a.countZ0Z_2\,
            ltout => OPEN,
            carryin => \a.count_1_cry_1\,
            carryout => \a.count_1_cry_2\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7004\,
            in2 => \_gnd_net_\,
            in3 => \N__6993\,
            lcout => \a.countZ0Z_3\,
            ltout => OPEN,
            carryin => \a.count_1_cry_2\,
            carryout => \a.count_1_cry_3\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7280\,
            in2 => \_gnd_net_\,
            in3 => \N__7269\,
            lcout => \a.countZ0Z_4\,
            ltout => OPEN,
            carryin => \a.count_1_cry_3\,
            carryout => \a.count_1_cry_4\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7265\,
            in2 => \_gnd_net_\,
            in3 => \N__7254\,
            lcout => \a.countZ0Z_5\,
            ltout => OPEN,
            carryin => \a.count_1_cry_4\,
            carryout => \a.count_1_cry_5\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7250\,
            in2 => \_gnd_net_\,
            in3 => \N__7239\,
            lcout => \a.countZ0Z_6\,
            ltout => OPEN,
            carryin => \a.count_1_cry_5\,
            carryout => \a.count_1_cry_6\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7235\,
            in2 => \_gnd_net_\,
            in3 => \N__7224\,
            lcout => \a.countZ0Z_7\,
            ltout => OPEN,
            carryin => \a.count_1_cry_6\,
            carryout => \a.count_1_cry_7\,
            clk => \N__14260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7214\,
            in2 => \_gnd_net_\,
            in3 => \N__7197\,
            lcout => \a.count_1_8\,
            ltout => OPEN,
            carryin => \a.count_1_cry_7\,
            carryout => \a.count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_9_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7193\,
            in2 => \_gnd_net_\,
            in3 => \N__7182\,
            lcout => \a.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \a.count_1_cry_9\,
            clk => \N__14254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_10_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7175\,
            in2 => \_gnd_net_\,
            in3 => \N__7158\,
            lcout => \a.count_1_10\,
            ltout => OPEN,
            carryin => \a.count_1_cry_9\,
            carryout => \a.count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_11_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7151\,
            in2 => \_gnd_net_\,
            in3 => \N__7134\,
            lcout => \a.count_1_11\,
            ltout => OPEN,
            carryin => \a.count_1_cry_10\,
            carryout => \a.count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_12_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7398\,
            in2 => \_gnd_net_\,
            in3 => \N__7380\,
            lcout => \a.count_1_12\,
            ltout => OPEN,
            carryin => \a.count_1_cry_11\,
            carryout => \a.count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_13_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7377\,
            in2 => \_gnd_net_\,
            in3 => \N__7359\,
            lcout => \a.count_1_13\,
            ltout => OPEN,
            carryin => \a.count_1_cry_12\,
            carryout => \a.count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNO_0_14_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7356\,
            in2 => \_gnd_net_\,
            in3 => \N__7338\,
            lcout => \a.count_1_14\,
            ltout => OPEN,
            carryin => \a.count_1_cry_13\,
            carryout => \a.count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_15_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7335\,
            in2 => \_gnd_net_\,
            in3 => \N__7323\,
            lcout => \a.countZ0Z_15\,
            ltout => OPEN,
            carryin => \a.count_1_cry_14\,
            carryout => \a.count_1_cry_15\,
            clk => \N__14254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_16_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7320\,
            in2 => \_gnd_net_\,
            in3 => \N__7308\,
            lcout => \a.countZ0Z_16\,
            ltout => OPEN,
            carryin => \a.count_1_cry_15\,
            carryout => \a.count_1_cry_16\,
            clk => \N__14254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_17_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7305\,
            in2 => \_gnd_net_\,
            in3 => \N__7293\,
            lcout => \a.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \a.count_1_cry_17\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_18_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7458\,
            in2 => \_gnd_net_\,
            in3 => \N__7290\,
            lcout => \a.countZ0Z_18\,
            ltout => OPEN,
            carryin => \a.count_1_cry_17\,
            carryout => \a.count_1_cry_18\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_19_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7416\,
            in2 => \_gnd_net_\,
            in3 => \N__7287\,
            lcout => \a.countZ0Z_19\,
            ltout => OPEN,
            carryin => \a.count_1_cry_18\,
            carryout => \a.count_1_cry_19\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_20_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7430\,
            in2 => \_gnd_net_\,
            in3 => \N__7284\,
            lcout => \a.countZ0Z_20\,
            ltout => OPEN,
            carryin => \a.count_1_cry_19\,
            carryout => \a.count_1_cry_20\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_21_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7445\,
            in2 => \_gnd_net_\,
            in3 => \N__7527\,
            lcout => \a.countZ0Z_21\,
            ltout => OPEN,
            carryin => \a.count_1_cry_20\,
            carryout => \a.count_1_cry_21\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_22_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7523\,
            in2 => \_gnd_net_\,
            in3 => \N__7509\,
            lcout => \a.countZ0Z_22\,
            ltout => OPEN,
            carryin => \a.count_1_cry_21\,
            carryout => \a.count_1_cry_22\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_23_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7506\,
            in2 => \_gnd_net_\,
            in3 => \N__7494\,
            lcout => \a.countZ0Z_23\,
            ltout => OPEN,
            carryin => \a.count_1_cry_22\,
            carryout => \a.count_1_cry_23\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_24_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7491\,
            in2 => \_gnd_net_\,
            in3 => \N__7479\,
            lcout => \a.countZ0Z_24\,
            ltout => OPEN,
            carryin => \a.count_1_cry_23\,
            carryout => \a.count_1_cry_24\,
            clk => \N__14247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_25_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7472\,
            in2 => \_gnd_net_\,
            in3 => \N__7476\,
            lcout => \a.countZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_1_c_RNO_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7562\,
            in1 => \N__7547\,
            in2 => \N__7581\,
            in3 => \N__7595\,
            lcout => decrement_time_0_prescaler10_1_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_0_c_RNO_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7614\,
            in1 => \N__7632\,
            in2 => \N__7677\,
            in3 => \N__7648\,
            lcout => decrement_time_0_prescaler10_0_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_RNIOGM61_18_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7457\,
            in1 => \N__7446\,
            in2 => \N__7431\,
            in3 => \N__7415\,
            lcout => \a.BUZZER3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_1_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7674\,
            in2 => \N__7653\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => prescaler_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_2_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7631\,
            in2 => \_gnd_net_\,
            in3 => \N__7617\,
            lcout => \prescalerZ0Z_2\,
            ltout => OPEN,
            carryin => prescaler_1_cry_1,
            carryout => prescaler_1_cry_2,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_3_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7613\,
            in2 => \_gnd_net_\,
            in3 => \N__7599\,
            lcout => \prescalerZ0Z_3\,
            ltout => OPEN,
            carryin => prescaler_1_cry_2,
            carryout => prescaler_1_cry_3,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_4_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7596\,
            in2 => \_gnd_net_\,
            in3 => \N__7584\,
            lcout => \prescalerZ0Z_4\,
            ltout => OPEN,
            carryin => prescaler_1_cry_3,
            carryout => prescaler_1_cry_4,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_5_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7580\,
            in2 => \_gnd_net_\,
            in3 => \N__7566\,
            lcout => \prescalerZ0Z_5\,
            ltout => OPEN,
            carryin => prescaler_1_cry_4,
            carryout => prescaler_1_cry_5,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_6_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7563\,
            in2 => \_gnd_net_\,
            in3 => \N__7551\,
            lcout => \prescalerZ0Z_6\,
            ltout => OPEN,
            carryin => prescaler_1_cry_5,
            carryout => prescaler_1_cry_6,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_7_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7548\,
            in2 => \_gnd_net_\,
            in3 => \N__7536\,
            lcout => \prescalerZ0Z_7\,
            ltout => OPEN,
            carryin => prescaler_1_cry_6,
            carryout => prescaler_1_cry_7,
            clk => \N__14233\,
            ce => \N__8055\,
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_7_THRU_LUT4_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7902\,
            in2 => \_gnd_net_\,
            in3 => \N__7533\,
            lcout => \prescaler_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_7,
            carryout => prescaler_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_9_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8468\,
            in2 => \_gnd_net_\,
            in3 => \N__7530\,
            lcout => \prescalerZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => prescaler_1_cry_9,
            clk => \N__14225\,
            ce => \N__8056\,
            sr => \_gnd_net_\
        );

    \prescaler_10_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8495\,
            in2 => \_gnd_net_\,
            in3 => \N__7704\,
            lcout => \prescalerZ0Z_10\,
            ltout => OPEN,
            carryin => prescaler_1_cry_9,
            carryout => prescaler_1_cry_10,
            clk => \N__14225\,
            ce => \N__8056\,
            sr => \_gnd_net_\
        );

    \prescaler_11_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8481\,
            in2 => \_gnd_net_\,
            in3 => \N__7701\,
            lcout => \prescalerZ0Z_11\,
            ltout => OPEN,
            carryin => prescaler_1_cry_10,
            carryout => prescaler_1_cry_11,
            clk => \N__14225\,
            ce => \N__8056\,
            sr => \_gnd_net_\
        );

    \prescaler_12_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8454\,
            in2 => \_gnd_net_\,
            in3 => \N__7698\,
            lcout => \prescalerZ0Z_12\,
            ltout => OPEN,
            carryin => prescaler_1_cry_11,
            carryout => prescaler_1_cry_12,
            clk => \N__14225\,
            ce => \N__8056\,
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_12_THRU_LUT4_0_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8202\,
            in2 => \_gnd_net_\,
            in3 => \N__7695\,
            lcout => \prescaler_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_12,
            carryout => prescaler_1_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_13_THRU_LUT4_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8163\,
            in2 => \_gnd_net_\,
            in3 => \N__7692\,
            lcout => \prescaler_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_13,
            carryout => prescaler_1_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_14_THRU_LUT4_0_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8127\,
            in2 => \_gnd_net_\,
            in3 => \N__7689\,
            lcout => \prescaler_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_14,
            carryout => prescaler_1_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_15_THRU_LUT4_0_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8094\,
            in2 => \_gnd_net_\,
            in3 => \N__7686\,
            lcout => \prescaler_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_15,
            carryout => prescaler_1_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_17_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8399\,
            in2 => \_gnd_net_\,
            in3 => \N__7683\,
            lcout => \prescalerZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => prescaler_1_cry_17,
            clk => \N__14219\,
            ce => \N__8057\,
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_17_THRU_LUT4_0_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7953\,
            in2 => \_gnd_net_\,
            in3 => \N__7680\,
            lcout => \prescaler_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_17,
            carryout => prescaler_1_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_19_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8385\,
            in2 => \_gnd_net_\,
            in3 => \N__7731\,
            lcout => \prescalerZ0Z_19\,
            ltout => OPEN,
            carryin => prescaler_1_cry_18,
            carryout => prescaler_1_cry_19,
            clk => \N__14219\,
            ce => \N__8057\,
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_19_THRU_LUT4_0_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8031\,
            in2 => \_gnd_net_\,
            in3 => \N__7728\,
            lcout => \prescaler_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_19,
            carryout => prescaler_1_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_20_THRU_LUT4_0_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8007\,
            in2 => \_gnd_net_\,
            in3 => \N__7725\,
            lcout => \prescaler_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_20,
            carryout => prescaler_1_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_21_THRU_LUT4_0_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7983\,
            in3 => \N__7722\,
            lcout => \prescaler_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_21,
            carryout => prescaler_1_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_22_THRU_LUT4_0_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7866\,
            in2 => \_gnd_net_\,
            in3 => \N__7719\,
            lcout => \prescaler_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_22,
            carryout => prescaler_1_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_23_THRU_LUT4_0_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7833\,
            in2 => \_gnd_net_\,
            in3 => \N__7716\,
            lcout => \prescaler_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_23,
            carryout => prescaler_1_cry_24,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_25_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8426\,
            in2 => \_gnd_net_\,
            in3 => \N__7713\,
            lcout => \prescalerZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => prescaler_1_cry_25,
            clk => \N__14215\,
            ce => \N__8058\,
            sr => \_gnd_net_\
        );

    \prescaler_1_cry_25_THRU_LUT4_0_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7791\,
            in2 => \_gnd_net_\,
            in3 => \N__7710\,
            lcout => \prescaler_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => prescaler_1_cry_25,
            carryout => prescaler_1_cry_26,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_27_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8412\,
            in2 => \_gnd_net_\,
            in3 => \N__7707\,
            lcout => \prescalerZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14215\,
            ce => \N__8058\,
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_4_c_RNO_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7891\,
            in1 => \N__7858\,
            in2 => \N__7829\,
            in3 => \N__7783\,
            lcout => decrement_time_0_prescaler10_4_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_8_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7901\,
            in1 => \N__7914\,
            in2 => \_gnd_net_\,
            in3 => \N__9944\,
            lcout => \prescalerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_23_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9941\,
            in1 => \N__7878\,
            in2 => \_gnd_net_\,
            in3 => \N__7859\,
            lcout => \prescalerZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_24_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7828\,
            in1 => \N__7845\,
            in2 => \_gnd_net_\,
            in3 => \N__9942\,
            lcout => \prescalerZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_26_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9943\,
            in1 => \N__7806\,
            in2 => \_gnd_net_\,
            in3 => \N__7784\,
            lcout => \prescalerZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_20_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7770\,
            in1 => \N__8027\,
            in2 => \_gnd_net_\,
            in3 => \N__9938\,
            lcout => \prescalerZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_21_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9939\,
            in1 => \N__7755\,
            in2 => \_gnd_net_\,
            in3 => \N__8003\,
            lcout => \prescalerZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \prescaler_22_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7743\,
            in1 => \N__7972\,
            in2 => \_gnd_net_\,
            in3 => \N__9940\,
            lcout => \prescalerZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14255\,
            ce => \N__8052\,
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_2_c_RNO_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8083\,
            in1 => \N__8119\,
            in2 => \N__8198\,
            in3 => \N__8155\,
            lcout => decrement_time_0_prescaler10_2_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescaler_13_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8197\,
            in1 => \N__8214\,
            in2 => \_gnd_net_\,
            in3 => \N__9915\,
            lcout => \prescalerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14248\,
            ce => \N__8054\,
            sr => \_gnd_net_\
        );

    \prescaler_14_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9916\,
            in1 => \N__8175\,
            in2 => \_gnd_net_\,
            in3 => \N__8156\,
            lcout => \prescalerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14248\,
            ce => \N__8054\,
            sr => \_gnd_net_\
        );

    \prescaler_15_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8120\,
            in1 => \N__8142\,
            in2 => \_gnd_net_\,
            in3 => \N__9917\,
            lcout => \prescalerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14248\,
            ce => \N__8054\,
            sr => \_gnd_net_\
        );

    \prescaler_16_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000010100"
        )
    port map (
            in0 => \N__9918\,
            in1 => \N__8106\,
            in2 => \N__8090\,
            in3 => \_gnd_net_\,
            lcout => \prescalerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14248\,
            ce => \N__8054\,
            sr => \_gnd_net_\
        );

    \prescaler_18_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7946\,
            in1 => \N__8070\,
            in2 => \_gnd_net_\,
            in3 => \N__9919\,
            lcout => \prescalerZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14248\,
            ce => \N__8054\,
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_3_c_RNO_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8023\,
            in1 => \N__7999\,
            in2 => \N__7979\,
            in3 => \N__7945\,
            lcout => decrement_time_0_prescaler10_3_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_0_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => decrement_time_0_prescaler10_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_1_c_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7923\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_0,
            carryout => decrement_time_0_prescaler10_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_2_c_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_1,
            carryout => decrement_time_0_prescaler10_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_3_c_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8238\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_2,
            carryout => decrement_time_0_prescaler10_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_4_c_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8229\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_3,
            carryout => decrement_time_0_prescaler10_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_5_c_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8442\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_4,
            carryout => decrement_time_0_prescaler10_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_6_c_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8373\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => decrement_time_0_prescaler10_5,
            carryout => decrement_time_0_prescaler10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_THRU_LUT4_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8217\,
            lcout => \decrement_time_0_prescaler10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_stored_e_0_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \mins_storedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14234\,
            ce => \N__10778\,
            sr => \_gnd_net_\
        );

    \mins_stored_e_0_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \mins_storedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14234\,
            ce => \N__10778\,
            sr => \_gnd_net_\
        );

    \mins_stored_e_0_2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13788\,
            lcout => \mins_storedZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14234\,
            ce => \N__10778\,
            sr => \_gnd_net_\
        );

    \d3.count_RNI1N275_12_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8727\,
            in1 => \N__8706\,
            in2 => \N__9699\,
            in3 => \N__8628\,
            lcout => d3_trans_up_1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_6_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13544\,
            in1 => \N__13885\,
            in2 => \N__13646\,
            in3 => \N__13756\,
            lcout => OPEN,
            ltout => \d1.mins27_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__12114\,
            in1 => \N__11124\,
            in2 => \N__8355\,
            in3 => \N__8508\,
            lcout => OPEN,
            ltout => \d1.g2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_0_o3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__10494\,
            in1 => \N__8322\,
            in2 => \N__8352\,
            in3 => \N__10024\,
            lcout => \d1.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ten_secs_2_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__10896\,
            in1 => \N__10589\,
            in2 => \N__12390\,
            in3 => \N__8747\,
            lcout => \ten_secsZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI5FPI2_3_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8349\,
            in1 => \N__8340\,
            in2 => \N__10945\,
            in3 => \N__8850\,
            lcout => \d1.g0_1_a5_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_11_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13757\,
            in1 => \N__13614\,
            in2 => \N__13897\,
            in3 => \N__13545\,
            lcout => \d1.g0_0_0_a4_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11084\,
            in2 => \_gnd_net_\,
            in3 => \N__9816\,
            lcout => \d1.gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIH1EH_7_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__8933\,
            in1 => \N__8315\,
            in2 => \N__8280\,
            in3 => \N__8875\,
            lcout => \d1.g1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIQ6A21_11_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8316\,
            in1 => \N__8276\,
            in2 => \N__8619\,
            in3 => \N__8849\,
            lcout => \d1.trans_up_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ten_secs_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10901\,
            in1 => \N__12429\,
            in2 => \_gnd_net_\,
            in3 => \N__8748\,
            lcout => \ten_secsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_2_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__11710\,
            in1 => \N__11284\,
            in2 => \N__12799\,
            in3 => \N__9237\,
            lcout => \d1.g2_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.sync_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8562\,
            lcout => \d3.syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_12_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12109\,
            in1 => \N__9258\,
            in2 => \N__12800\,
            in3 => \N__12356\,
            lcout => OPEN,
            ltout => \d1.g2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_0_4_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8550\,
            in2 => \N__8502\,
            in3 => \N__11285\,
            lcout => \d1.g2_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_5_c_RNO_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8499\,
            in1 => \N__8480\,
            in2 => \N__8469\,
            in3 => \N__8453\,
            lcout => decrement_time_0_prescaler10_5_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \decrement_time_0_prescaler10_6_c_RNO_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__8411\,
            in2 => \N__8400\,
            in3 => \N__8384\,
            lcout => decrement_time_0_prescaler10_6_and,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_15_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11493\,
            in1 => \N__11634\,
            in2 => \N__11712\,
            in3 => \N__11440\,
            lcout => OPEN,
            ltout => \d1.g2_7_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_11_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__11237\,
            in1 => \N__11180\,
            in2 => \N__8358\,
            in3 => \N__11903\,
            lcout => \d1.g2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNID2KP_9_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__8612\,
            in1 => \N__8903\,
            in2 => \N__9076\,
            in3 => \N__8960\,
            lcout => \d1.g1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIVLG6B_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__11541\,
            in1 => \N__10161\,
            in2 => \N__10188\,
            in3 => \N__10124\,
            lcout => \d1.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.sync_0_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8580\,
            lcout => \d3.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_5_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11492\,
            in1 => \N__11622\,
            in2 => \N__11711\,
            in3 => \N__11434\,
            lcout => \d1.g2_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8541\,
            lcout => d2_sync_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_1_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11626\,
            in2 => \_gnd_net_\,
            in3 => \N__11439\,
            lcout => d2_count_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14207\,
            ce => 'H',
            sr => \N__10290\
        );

    \d2.count_0_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11438\,
            lcout => d2_count_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14207\,
            ce => 'H',
            sr => \N__10290\
        );

    \d4.sync_1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13311\,
            lcout => \d4.syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.sync_1_RNIQPEK_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8721\,
            in2 => \_gnd_net_\,
            in3 => \N__8795\,
            lcout => \d4.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9362\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9337\,
            lcout => \d4.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14256\,
            ce => 'H',
            sr => \N__9619\
        );

    \d4.count_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9361\,
            lcout => \d4.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14256\,
            ce => 'H',
            sr => \N__9619\
        );

    \d1.g2_9_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13780\,
            in1 => \N__13671\,
            in2 => \N__13547\,
            in3 => \N__13898\,
            lcout => OPEN,
            ltout => \d1.g2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_0_3_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__11882\,
            in1 => \N__11238\,
            in2 => \N__8670\,
            in3 => \N__11181\,
            lcout => \d1.g2_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.ten_secs_1_sqmuxa_0_x1_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12494\,
            in1 => \N__12449\,
            in2 => \N__10607\,
            in3 => \N__11881\,
            lcout => OPEN,
            ltout => \d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.ten_secs_1_sqmuxa_0_ns_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8667\,
            in3 => \N__12759\,
            lcout => \d1.ten_secs_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a.count_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8655\,
            lcout => \a.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_RNI5PSB_10_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9467\,
            in1 => \N__9452\,
            in2 => \N__9438\,
            in3 => \N__9482\,
            lcout => \d4.trans_up_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_RNIS9LE1_10_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__9738\,
            in1 => \N__9580\,
            in2 => \N__9720\,
            in3 => \N__9603\,
            lcout => \d3.trans_up_1_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9605\,
            in1 => \_gnd_net_\,
            in2 => \N__9587\,
            in3 => \_gnd_net_\,
            lcout => \d3.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14240\,
            ce => 'H',
            sr => \N__9958\
        );

    \d3.count_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9604\,
            lcout => \d3.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14240\,
            ce => 'H',
            sr => \N__9958\
        );

    \d4.count_RNICSOB_16_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9653\,
            in1 => \N__9314\,
            in2 => \N__9636\,
            in3 => \N__9338\,
            lcout => \d4.trans_up_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_RNIE50C_3_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9284\,
            in1 => \N__9269\,
            in2 => \N__9501\,
            in3 => \N__9299\,
            lcout => \d4.trans_up_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_RNIMDFN1_6_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9770\,
            in1 => \N__9785\,
            in2 => \N__9756\,
            in3 => \N__9800\,
            lcout => \d3.trans_up_1_15_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.sync_1_RNIHL7Q_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__9386\,
            in1 => \N__8720\,
            in2 => \N__9672\,
            in3 => \N__8792\,
            lcout => \d4.trans_up_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_RNI6TEN1_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__9551\,
            in2 => \N__9522\,
            in3 => \N__9566\,
            lcout => \d3.trans_up_1_15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.state_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8763\,
            in2 => \_gnd_net_\,
            in3 => \N__8794\,
            lcout => d4_state,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_RNIFDLK_11_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9419\,
            in1 => \N__9366\,
            in2 => \N__9405\,
            in3 => \N__8700\,
            lcout => OPEN,
            ltout => \d4.trans_up_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_RNIQ4M62_11_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8691\,
            in1 => \N__8685\,
            in2 => \N__8679\,
            in3 => \N__8676\,
            lcout => d4_trans_up_1,
            ltout => \d4_trans_up_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_1_sqmuxa_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__8793\,
            in1 => \_gnd_net_\,
            in2 => \N__8808\,
            in3 => \N__9865\,
            lcout => \d1.state_1_sqmuxaZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ten_secs_RNO_0_1_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8743\,
            lcout => OPEN,
            ltout => \ten_secs_r_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ten_secs_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__10902\,
            in1 => \N__12490\,
            in2 => \N__8805\,
            in3 => \N__10825\,
            lcout => \ten_secsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_RNIEJS51_16_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10666\,
            in1 => \N__10649\,
            in2 => \N__9837\,
            in3 => \N__10631\,
            lcout => \d3.trans_up_1_14_2\,
            ltout => \d3.trans_up_1_14_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.state_RNI7N9P6_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12576\,
            in1 => \N__12609\,
            in2 => \N__8802\,
            in3 => \N__11083\,
            lcout => s_cancel,
            ltout => \s_cancel_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.alarm_on_0_sqmuxa_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12770\,
            in2 => \N__8799\,
            in3 => \N__11886\,
            lcout => alarm_on_0_sqmuxa,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.mins_stored_0_sqmuxa_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11888\,
            in1 => \N__8796\,
            in2 => \N__12796\,
            in3 => \N__8762\,
            lcout => mins_stored_0_sqmuxa,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.secs_0_sqmuxa_ns_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10095\,
            in2 => \_gnd_net_\,
            in3 => \N__9911\,
            lcout => secs_0_sqmuxa,
            ltout => \secs_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.un1_state_9_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000001000000"
        )
    port map (
            in0 => \N__11887\,
            in1 => \N__12789\,
            in2 => \N__8751\,
            in3 => \N__9869\,
            lcout => un1_state_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__11082\,
            in1 => \N__9812\,
            in2 => \N__9012\,
            in3 => \N__10023\,
            lcout => ten_secs_1_sqmuxa,
            ltout => \ten_secs_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_0_0_1_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100001110"
        )
    port map (
            in0 => \N__9000\,
            in1 => \N__8994\,
            in2 => \N__8985\,
            in3 => \N__13631\,
            lcout => OPEN,
            ltout => \d1.g0_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNI7SNV11_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000001111"
        )
    port map (
            in0 => \N__8982\,
            in1 => \N__10062\,
            in2 => \N__8973\,
            in3 => \N__13543\,
            lcout => OPEN,
            ltout => \d1.un1_mins_4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_1_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__8970\,
            in1 => \N__11115\,
            in2 => \N__8964\,
            in3 => \N__9870\,
            lcout => \minsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14221\,
            ce => 'H',
            sr => \N__11564\
        );

    \d1.count_RNIP9EH_7_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8961\,
            in1 => \N__8934\,
            in2 => \N__8907\,
            in3 => \N__8877\,
            lcout => \d1.trans_up_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_8_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__10194\,
            in1 => \N__8838\,
            in2 => \N__10826\,
            in3 => \N__11505\,
            lcout => \d1.un1_mins_1_sqmuxa_0\,
            ltout => \d1.un1_mins_1_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNID20IK_3_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__10911\,
            in1 => \N__9198\,
            in2 => \N__8832\,
            in3 => \N__10163\,
            lcout => OPEN,
            ltout => \d1.un1_mins_3_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI7SNV11_3_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100001000"
        )
    port map (
            in0 => \N__13632\,
            in1 => \N__13511\,
            in2 => \N__8829\,
            in3 => \N__8826\,
            lcout => OPEN,
            ltout => \d1.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_2_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__8820\,
            in1 => \N__13772\,
            in2 => \N__8811\,
            in3 => \N__10892\,
            lcout => \minsZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14216\,
            ce => 'H',
            sr => \N__11551\
        );

    \d1.count_RNI0GQ42_7_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__9213\,
            in1 => \N__10041\,
            in2 => \N__9207\,
            in3 => \N__9152\,
            lcout => \d1.g1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIH6847_16_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9192\,
            in1 => \N__9180\,
            in2 => \N__11520\,
            in3 => \N__10153\,
            lcout => \d1.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI1SGU2_3_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9171\,
            in1 => \N__10946\,
            in2 => \N__9153\,
            in3 => \N__9119\,
            lcout => \d1.trans_up_1_0\,
            ltout => \d1.trans_up_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNISBML3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__9080\,
            in1 => \N__12785\,
            in2 => \N__9108\,
            in3 => \N__11904\,
            lcout => \d1.g0_2_0_o2_2\,
            ltout => \d1.g0_2_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIA71EK_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000110111"
        )
    port map (
            in0 => \N__10154\,
            in1 => \N__10061\,
            in2 => \N__9105\,
            in3 => \N__13503\,
            lcout => OPEN,
            ltout => \d1.N_19_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__9102\,
            in1 => \N__9090\,
            in2 => \N__9084\,
            in3 => \N__10897\,
            lcout => \minsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_2_0_a4_2_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13765\,
            in1 => \N__13651\,
            in2 => \N__13535\,
            in3 => \N__13892\,
            lcout => \d1.g0_2_0_a4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNI4LMC_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13650\,
            in1 => \N__13499\,
            in2 => \N__9081\,
            in3 => \N__13764\,
            lcout => \d1.g2_i_a5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_RNIP8VS_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12246\,
            in1 => \N__12017\,
            in2 => \N__11958\,
            in3 => \N__11752\,
            lcout => \d2.g0_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_6_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__11751\,
            in1 => \N__11945\,
            in2 => \N__12032\,
            in3 => \N__12245\,
            lcout => \d1.g2_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNI1DIH_13_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11427\,
            in1 => \N__12151\,
            in2 => \N__12177\,
            in3 => \N__11479\,
            lcout => OPEN,
            ltout => \d2.g0_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIJ0PB1_8_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11165\,
            in1 => \N__11306\,
            in2 => \N__9249\,
            in3 => \N__11221\,
            lcout => OPEN,
            ltout => \d2.g0_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIK9TB3_10_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12258\,
            in1 => \N__9246\,
            in2 => \N__9240\,
            in3 => \N__9228\,
            lcout => s_dn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__12018\,
            in1 => \N__11388\,
            in2 => \N__9222\,
            in3 => \N__11949\,
            lcout => d2_state,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNI3QT21_4_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11426\,
            in1 => \N__11480\,
            in2 => \N__11230\,
            in3 => \N__11164\,
            lcout => d2_trans_up_1_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_4_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11478\,
            in1 => \N__11608\,
            in2 => \N__11761\,
            in3 => \N__11425\,
            lcout => \d1.g2_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIS7IH_11_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12135\,
            in1 => \N__11680\,
            in2 => \N__12198\,
            in3 => \N__11620\,
            lcout => \d2.g0_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNO_0_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11621\,
            in1 => \N__12337\,
            in2 => \N__11697\,
            in3 => \N__12248\,
            lcout => \d2.trans_up_1_14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_7_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11217\,
            in1 => \N__11163\,
            in2 => \N__12348\,
            in3 => \N__12242\,
            lcout => OPEN,
            ltout => \d1.g2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_0_3_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__12025\,
            in1 => \_gnd_net_\,
            in2 => \N__9372\,
            in3 => \N__12790\,
            lcout => \d1.g2_i_a5_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_0_a4_7_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11335\,
            in1 => \N__13781\,
            in2 => \N__13546\,
            in3 => \N__11759\,
            lcout => OPEN,
            ltout => \d1.g0_1_0_a4Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_0_a4_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11775\,
            in1 => \N__12113\,
            in2 => \N__9369\,
            in3 => \N__11286\,
            lcout => mins_0_sqmuxa,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.un3_count_cry_1_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9360\,
            in2 => \N__9339\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \d4.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d4.count_2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9315\,
            in2 => \_gnd_net_\,
            in3 => \N__9303\,
            lcout => \d4.countZ0Z_2\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_1\,
            carryout => \d4.un3_count_cry_2\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9300\,
            in2 => \_gnd_net_\,
            in3 => \N__9288\,
            lcout => \d4.countZ0Z_3\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_2\,
            carryout => \d4.un3_count_cry_3\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_4_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9285\,
            in2 => \_gnd_net_\,
            in3 => \N__9273\,
            lcout => \d4.countZ0Z_4\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_3\,
            carryout => \d4.un3_count_cry_4\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9270\,
            in2 => \_gnd_net_\,
            in3 => \N__9504\,
            lcout => \d4.countZ0Z_5\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_4\,
            carryout => \d4.un3_count_cry_5\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_6_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9500\,
            in2 => \_gnd_net_\,
            in3 => \N__9486\,
            lcout => \d4.countZ0Z_6\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_5\,
            carryout => \d4.un3_count_cry_6\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_7_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9483\,
            in2 => \_gnd_net_\,
            in3 => \N__9471\,
            lcout => \d4.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_6\,
            carryout => \d4.un3_count_cry_7\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9468\,
            in2 => \_gnd_net_\,
            in3 => \N__9456\,
            lcout => \d4.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_7\,
            carryout => \d4.un3_count_cry_8\,
            clk => \N__14241\,
            ce => 'H',
            sr => \N__9620\
        );

    \d4.count_9_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9453\,
            in2 => \_gnd_net_\,
            in3 => \N__9441\,
            lcout => \d4.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \d4.un3_count_cry_9\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_10_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9437\,
            in2 => \_gnd_net_\,
            in3 => \N__9423\,
            lcout => \d4.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_9\,
            carryout => \d4.un3_count_cry_10\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_11_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9420\,
            in2 => \_gnd_net_\,
            in3 => \N__9408\,
            lcout => \d4.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_10\,
            carryout => \d4.un3_count_cry_11\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_12_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9404\,
            in2 => \_gnd_net_\,
            in3 => \N__9390\,
            lcout => \d4.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_11\,
            carryout => \d4.un3_count_cry_12\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_13_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9387\,
            in2 => \_gnd_net_\,
            in3 => \N__9375\,
            lcout => \d4.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_12\,
            carryout => \d4.un3_count_cry_13\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_14_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9671\,
            in2 => \_gnd_net_\,
            in3 => \N__9657\,
            lcout => \d4.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_13\,
            carryout => \d4.un3_count_cry_14\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_15_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9654\,
            in2 => \_gnd_net_\,
            in3 => \N__9642\,
            lcout => \d4.countZ0Z_15\,
            ltout => OPEN,
            carryin => \d4.un3_count_cry_14\,
            carryout => \d4.un3_count_cry_15\,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d4.count_16_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9635\,
            in2 => \_gnd_net_\,
            in3 => \N__9639\,
            lcout => \d4.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14236\,
            ce => 'H',
            sr => \N__9621\
        );

    \d3.un3_count_cry_1_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9606\,
            in2 => \N__9588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \d3.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9567\,
            in2 => \_gnd_net_\,
            in3 => \N__9555\,
            lcout => \d3.countZ0Z_2\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_1\,
            carryout => \d3.un3_count_cry_2\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_3_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9552\,
            in2 => \_gnd_net_\,
            in3 => \N__9540\,
            lcout => \d3.countZ0Z_3\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_2\,
            carryout => \d3.un3_count_cry_3\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9537\,
            in2 => \_gnd_net_\,
            in3 => \N__9525\,
            lcout => \d3.countZ0Z_4\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_3\,
            carryout => \d3.un3_count_cry_4\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9521\,
            in2 => \_gnd_net_\,
            in3 => \N__9507\,
            lcout => \d3.countZ0Z_5\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_4\,
            carryout => \d3.un3_count_cry_5\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_6_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9801\,
            in2 => \_gnd_net_\,
            in3 => \N__9789\,
            lcout => \d3.countZ0Z_6\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_5\,
            carryout => \d3.un3_count_cry_6\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9786\,
            in2 => \_gnd_net_\,
            in3 => \N__9774\,
            lcout => \d3.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_6\,
            carryout => \d3.un3_count_cry_7\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9771\,
            in2 => \_gnd_net_\,
            in3 => \N__9759\,
            lcout => \d3.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_7\,
            carryout => \d3.un3_count_cry_8\,
            clk => \N__14228\,
            ce => 'H',
            sr => \N__9959\
        );

    \d3.count_9_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9755\,
            in2 => \_gnd_net_\,
            in3 => \N__9741\,
            lcout => \d3.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \d3.un3_count_cry_9\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_10_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9737\,
            in2 => \_gnd_net_\,
            in3 => \N__9723\,
            lcout => \d3.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_9\,
            carryout => \d3.un3_count_cry_10\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_11_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9716\,
            in2 => \_gnd_net_\,
            in3 => \N__9702\,
            lcout => \d3.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_10\,
            carryout => \d3.un3_count_cry_11\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9695\,
            in2 => \_gnd_net_\,
            in3 => \N__9681\,
            lcout => \d3.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_11\,
            carryout => \d3.un3_count_cry_12\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_13_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9836\,
            in2 => \_gnd_net_\,
            in3 => \N__9678\,
            lcout => \d3.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_12\,
            carryout => \d3.un3_count_cry_13\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_14_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10632\,
            in2 => \_gnd_net_\,
            in3 => \N__9675\,
            lcout => \d3.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_13\,
            carryout => \d3.un3_count_cry_14\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_15_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10650\,
            in2 => \_gnd_net_\,
            in3 => \N__9966\,
            lcout => \d3.countZ0Z_15\,
            ltout => OPEN,
            carryin => \d3.un3_count_cry_14\,
            carryout => \d3.un3_count_cry_15\,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d3.count_16_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10668\,
            in2 => \_gnd_net_\,
            in3 => \N__9963\,
            lcout => \d3.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14222\,
            ce => 'H',
            sr => \N__9960\
        );

    \d1.un1_state_7_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000000000"
        )
    port map (
            in0 => \N__9868\,
            in1 => \N__11891\,
            in2 => \N__12801\,
            in3 => \N__9945\,
            lcout => un1_state_7_0,
            ltout => \un1_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101000000000"
        )
    port map (
            in0 => \N__10442\,
            in1 => \N__10351\,
            in2 => \N__9882\,
            in3 => \N__9876\,
            lcout => \secsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.un1_alarm_on_0_sqmuxa_0_i_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__12795\,
            in1 => \N__9866\,
            in2 => \_gnd_net_\,
            in3 => \N__11889\,
            lcout => un1_alarm_on_0_sqmuxa_0_i,
            ltout => \un1_alarm_on_0_sqmuxa_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_RNO_0_1_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10534\,
            in2 => \N__9879\,
            in3 => \N__10025\,
            lcout => \N_120_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_0_sqmuxa_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13542\,
            in1 => \N__13866\,
            in2 => \N__13634\,
            in3 => \N__13776\,
            lcout => \d1.state_0_sqmuxaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_2_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111111111"
        )
    port map (
            in0 => \N__11890\,
            in1 => \N__12791\,
            in2 => \_gnd_net_\,
            in3 => \N__9867\,
            lcout => un1_alarm_on_0_sqmuxa_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.state_RNI607I1_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12567\,
            in1 => \N__9832\,
            in2 => \N__12617\,
            in3 => \N__10614\,
            lcout => d3_g0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.secs_0_sqmuxa_x1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10469\,
            in1 => \N__10435\,
            in2 => \N__10399\,
            in3 => \N__10350\,
            lcout => \d1.secs_0_sqmuxa_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.mins_16_1_3_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011110001011"
        )
    port map (
            in0 => \N__13849\,
            in1 => \N__10878\,
            in2 => \N__10086\,
            in3 => \N__10060\,
            lcout => \d1.mins_16_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__10358\,
            in1 => \N__9999\,
            in2 => \_gnd_net_\,
            in3 => \N__9976\,
            lcout => \secsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIC9AJK_16_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__13510\,
            in1 => \N__10068\,
            in2 => \N__12522\,
            in3 => \N__10059\,
            lcout => \d1.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_10_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13487\,
            in1 => \N__13848\,
            in2 => \N__13680\,
            in3 => \N__13755\,
            lcout => \d1.g0_0_0_a4_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_RNO_0_2_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__10473\,
            in1 => \N__10440\,
            in2 => \N__10001\,
            in3 => \N__10356\,
            lcout => OPEN,
            ltout => \secs_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_2_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__9978\,
            in2 => \N__10032\,
            in3 => \N__10029\,
            lcout => \secsZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_RNO_0_3_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__10474\,
            in1 => \N__10441\,
            in2 => \N__10002\,
            in3 => \N__10357\,
            lcout => OPEN,
            ltout => \un1_secs_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_3_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010010110"
        )
    port map (
            in0 => \N__10398\,
            in1 => \N__10000\,
            in2 => \N__9981\,
            in3 => \N__9977\,
            lcout => \secsZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIGDI57_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10217\,
            in1 => \N__10101\,
            in2 => \N__10206\,
            in3 => \N__11370\,
            lcout => \d1.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_9_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13748\,
            in1 => \N__13488\,
            in2 => \N__13681\,
            in3 => \N__13850\,
            lcout => \d1.mins27_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_0_1_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13841\,
            in2 => \_gnd_net_\,
            in3 => \N__13747\,
            lcout => OPEN,
            ltout => \d1.g0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_10_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011111111"
        )
    port map (
            in0 => \N__13670\,
            in1 => \N__13489\,
            in2 => \N__10197\,
            in3 => \N__11269\,
            lcout => \d1.g2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIINS67_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10187\,
            in1 => \N__10162\,
            in2 => \_gnd_net_\,
            in3 => \N__10125\,
            lcout => \d1.mins_2_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_0_6_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11696\,
            in1 => \N__10113\,
            in2 => \N__11985\,
            in3 => \N__11900\,
            lcout => OPEN,
            ltout => \d1.g2_i_a5_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_0_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__11349\,
            in1 => \N__11313\,
            in2 => \N__10104\,
            in3 => \N__12054\,
            lcout => \d1.g2_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_2_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11899\,
            lcout => \d1.g2_i_a5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.un3_count_cry_1_c_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11448\,
            in2 => \N__11643\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \d2.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_2_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11694\,
            in2 => \_gnd_net_\,
            in3 => \N__10248\,
            lcout => d2_count_2,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_1\,
            carryout => \d2.un3_count_cry_2\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_3_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12247\,
            in2 => \_gnd_net_\,
            in3 => \N__10245\,
            lcout => d2_count_3,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_2\,
            carryout => \d2.un3_count_cry_3\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_4_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11488\,
            in2 => \_gnd_net_\,
            in3 => \N__10242\,
            lcout => d2_count_4,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_3\,
            carryout => \d2.un3_count_cry_4\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_5_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11172\,
            in2 => \_gnd_net_\,
            in3 => \N__10239\,
            lcout => d2_count_5,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_4\,
            carryout => \d2.un3_count_cry_5\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_6_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11228\,
            in2 => \_gnd_net_\,
            in3 => \N__10236\,
            lcout => d2_count_6,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_5\,
            carryout => \d2.un3_count_cry_6\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_7_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12273\,
            in2 => \_gnd_net_\,
            in3 => \N__10233\,
            lcout => \d2.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_6\,
            carryout => \d2.un3_count_cry_7\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_8_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11307\,
            in2 => \_gnd_net_\,
            in3 => \N__10230\,
            lcout => \d2.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_7\,
            carryout => \d2.un3_count_cry_8\,
            clk => \N__14205\,
            ce => 'H',
            sr => \N__10289\
        );

    \d2.count_9_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12372\,
            in2 => \_gnd_net_\,
            in3 => \N__10227\,
            lcout => \d2.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \d2.un3_count_cry_9\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_10_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12292\,
            in2 => \_gnd_net_\,
            in3 => \N__10224\,
            lcout => \d2.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_9\,
            carryout => \d2.un3_count_cry_10\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_11_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12134\,
            in2 => \_gnd_net_\,
            in3 => \N__10308\,
            lcout => \d2.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_10\,
            carryout => \d2.un3_count_cry_11\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_12_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12197\,
            in2 => \_gnd_net_\,
            in3 => \N__10305\,
            lcout => \d2.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_11\,
            carryout => \d2.un3_count_cry_12\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_13_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12176\,
            in2 => \_gnd_net_\,
            in3 => \N__10302\,
            lcout => \d2.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_12\,
            carryout => \d2.un3_count_cry_13\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_14_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12155\,
            in2 => \_gnd_net_\,
            in3 => \N__10299\,
            lcout => \d2.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_13\,
            carryout => \d2.un3_count_cry_14\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_15_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11760\,
            in2 => \_gnd_net_\,
            in3 => \N__10296\,
            lcout => d2_count_15,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_14\,
            carryout => \d2.un3_count_cry_15\,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \d2.count_16_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12341\,
            in2 => \_gnd_net_\,
            in3 => \N__10293\,
            lcout => d2_count_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14204\,
            ce => 'H',
            sr => \N__10288\
        );

    \state_e_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10731\,
            in1 => \N__10323\,
            in2 => \_gnd_net_\,
            in3 => \N__10549\,
            lcout => \stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14223\,
            ce => \N__10275\,
            sr => \_gnd_net_\
        );

    \state_sbtinv_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10254\,
            lcout => un1_state_0_sqmuxa_1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.un1_state_0_sqmuxa_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__10719\,
            in1 => \N__10263\,
            in2 => \N__10545\,
            in3 => \N__10710\,
            lcout => un1_state_0_sqmuxa_1_0,
            ltout => \un1_state_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10782\,
            in3 => \N__12716\,
            lcout => \stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14218\,
            ce => 'H',
            sr => \N__10779\
        );

    \d1.state_0_sqmuxa_2_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10608\,
            in1 => \N__12495\,
            in2 => \N__10743\,
            in3 => \N__12450\,
            lcout => \d1.state_0_sqmuxaZ0Z_2\,
            ltout => \d1.state_0_sqmuxaZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_0_sqmuxa_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10319\,
            in2 => \N__10722\,
            in3 => \N__10530\,
            lcout => state_0_sqmuxa,
            ltout => \state_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alarm_on_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10682\,
            in2 => \N__10713\,
            in3 => \N__10709\,
            lcout => \alarm_onZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.count_RNI4GDS_16_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10667\,
            in1 => \N__10648\,
            in2 => \_gnd_net_\,
            in3 => \N__10630\,
            lcout => \d3.count_RNI4GDSZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.un1_state_3_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11860\,
            in2 => \_gnd_net_\,
            in3 => \N__12684\,
            lcout => un1_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_0_2_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__12505\,
            in2 => \N__10544\,
            in3 => \N__12451\,
            lcout => \d1.g0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secs_RNIUG5J_3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10478\,
            in1 => \N__10436\,
            in2 => \N__10400\,
            in3 => \N__10352\,
            lcout => decrement_time_0_secs9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_3_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11229\,
            in1 => \N__11173\,
            in2 => \N__12357\,
            in3 => \N__12249\,
            lcout => OPEN,
            ltout => \d1.g2_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__12047\,
            in1 => \N__11981\,
            in2 => \N__11127\,
            in3 => \N__11861\,
            lcout => \d1.g2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_13_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12749\,
            lcout => \d1.N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.state_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__12618\,
            in1 => \N__12575\,
            in2 => \N__11106\,
            in3 => \N__11091\,
            lcout => \d3.stateZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI2PCE_1_3_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11061\,
            in1 => \N__11034\,
            in2 => \N__11007\,
            in3 => \N__10974\,
            lcout => OPEN,
            ltout => \d1.g1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIUT4M1_3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10950\,
            in1 => \N__11901\,
            in2 => \N__10914\,
            in3 => \N__12748\,
            lcout => \d1.g1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNIKMMMV_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__10845\,
            in2 => \N__10839\,
            in3 => \N__10830\,
            lcout => OPEN,
            ltout => \d1.g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mins_3_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001010000010001"
        )
    port map (
            in0 => \N__10803\,
            in1 => \N__10797\,
            in2 => \N__10791\,
            in3 => \N__10788\,
            lcout => \minsZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14206\,
            ce => 'H',
            sr => \N__11568\
        );

    \d1.g0_1_a5_0_11_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12774\,
            in1 => \N__13862\,
            in2 => \N__13548\,
            in3 => \N__11898\,
            lcout => \d1.g0_1_a5_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_14_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12100\,
            in1 => \N__12204\,
            in2 => \N__12797\,
            in3 => \N__12352\,
            lcout => \d1.g2_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_8_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11484\,
            in1 => \N__11638\,
            in2 => \N__11766\,
            in3 => \N__11447\,
            lcout => \d1.g2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNID7FT1_15_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11343\,
            in1 => \N__11765\,
            in2 => \N__12102\,
            in3 => \N__11270\,
            lcout => \d2.trans_up_1_15\,
            ltout => \d2.trans_up_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIK9TB3_1_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11919\,
            in1 => \N__11639\,
            in2 => \N__11373\,
            in3 => \N__11695\,
            lcout => s_dn_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_0_7_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11364\,
            in1 => \N__12101\,
            in2 => \N__11358\,
            in3 => \N__11271\,
            lcout => \d1.g2_i_a5_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIQ9VS_16_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12244\,
            in1 => \N__11973\,
            in2 => \N__12046\,
            in3 => \N__12327\,
            lcout => d2_g0_3,
            ltout => \d2_g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_1_7_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12096\,
            in1 => \N__11342\,
            in2 => \N__11316\,
            in3 => \N__11272\,
            lcout => \d1.g2_i_a5_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNITE8Q_10_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12370\,
            in1 => \N__11299\,
            in2 => \N__12293\,
            in3 => \N__12271\,
            lcout => d2_trans_up_1_15_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNICOIH_10_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12371\,
            in1 => \N__12326\,
            in2 => \N__12294\,
            in3 => \N__12272\,
            lcout => \d2.g0_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_16_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__11972\,
            in1 => \N__11753\,
            in2 => \N__12045\,
            in3 => \N__12243\,
            lcout => \d1.g2_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNI237_11_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12193\,
            in1 => \N__12175\,
            in2 => \N__12156\,
            in3 => \N__12130\,
            lcout => d2_trans_up_1_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_1_6_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13550\,
            in1 => \N__12624\,
            in2 => \N__13682\,
            in3 => \N__11864\,
            lcout => \d1.g2_i_a5_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_RNIMV5K_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__12048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11980\,
            lcout => \d2.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_0_a4_4_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__13867\,
            in1 => \N__11684\,
            in2 => \N__13679\,
            in3 => \N__11628\,
            lcout => OPEN,
            ltout => \d1.g0_1_0_a4Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_0_a4_8_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11918\,
            in1 => \N__12731\,
            in2 => \N__11907\,
            in3 => \N__11863\,
            lcout => \d1.g0_1_0_a4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIOJGH_15_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11747\,
            in1 => \N__11685\,
            in2 => \_gnd_net_\,
            in3 => \N__11627\,
            lcout => OPEN,
            ltout => \d2_g0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g2_i_a5_1_3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12732\,
            in2 => \N__12627\,
            in3 => \N__13789\,
            lcout => \d1.g2_i_a5_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__13984\,
            in1 => \N__13074\,
            in2 => \N__14043\,
            in3 => \N__12813\,
            lcout => \display2.prescalerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNI3D3L_23_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12824\,
            in1 => \N__12848\,
            in2 => \N__13017\,
            in3 => \N__12872\,
            lcout => \display2.prescaler8_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_6_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__12837\,
            in1 => \N__14038\,
            in2 => \N__13083\,
            in3 => \N__13983\,
            lcout => \display2.prescalerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_4_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__12861\,
            in1 => \N__14037\,
            in2 => \N__13082\,
            in3 => \N__13982\,
            lcout => \display2.prescalerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d3.state_RNIOCAC_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12610\,
            in2 => \_gnd_net_\,
            in3 => \N__12568\,
            lcout => \d3.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.g0_1_0_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13675\,
            in2 => \_gnd_net_\,
            in3 => \N__13790\,
            lcout => \d1.g0_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.BNC1_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12506\,
            in2 => \_gnd_net_\,
            in3 => \N__12452\,
            lcout => \BNC1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_2_cry_1_c_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13101\,
            in2 => \N__13206\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \display2.prescaler_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_2_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12918\,
            in2 => \_gnd_net_\,
            in3 => \N__12879\,
            lcout => \display2.prescalerZ0Z_2\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_1\,
            carryout => \display2.prescaler_2_cry_2\,
            clk => \N__14242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_3_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12945\,
            in2 => \_gnd_net_\,
            in3 => \N__12876\,
            lcout => \display2.prescalerZ0Z_3\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_2\,
            carryout => \display2.prescaler_2_cry_3\,
            clk => \N__14242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_4_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12873\,
            in2 => \_gnd_net_\,
            in3 => \N__12855\,
            lcout => \display2.prescaler_2_4\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_3\,
            carryout => \display2.prescaler_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_5_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12957\,
            in2 => \_gnd_net_\,
            in3 => \N__12852\,
            lcout => \display2.prescalerZ0Z_5\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_4\,
            carryout => \display2.prescaler_2_cry_5\,
            clk => \N__14242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_6_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12849\,
            in2 => \_gnd_net_\,
            in3 => \N__12831\,
            lcout => \display2.prescaler_2_6\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_5\,
            carryout => \display2.prescaler_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_7_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12932\,
            in2 => \_gnd_net_\,
            in3 => \N__12828\,
            lcout => \display2.prescalerZ0Z_7\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_6\,
            carryout => \display2.prescaler_2_cry_7\,
            clk => \N__14242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_8_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12825\,
            in2 => \_gnd_net_\,
            in3 => \N__12807\,
            lcout => \display2.prescaler_2_8\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_7\,
            carryout => \display2.prescaler_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_9_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13173\,
            in2 => \_gnd_net_\,
            in3 => \N__12804\,
            lcout => \display2.prescaler_2_9\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \display2.prescaler_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_10_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13269\,
            in2 => \_gnd_net_\,
            in3 => \N__12906\,
            lcout => \display2.prescalerZ0Z_10\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_9\,
            carryout => \display2.prescaler_2_cry_10\,
            clk => \N__14237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_11_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13239\,
            in2 => \_gnd_net_\,
            in3 => \N__12903\,
            lcout => \display2.prescalerZ0Z_11\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_10\,
            carryout => \display2.prescaler_2_cry_11\,
            clk => \N__14237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_12_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13283\,
            in2 => \_gnd_net_\,
            in3 => \N__12900\,
            lcout => \display2.prescalerZ0Z_12\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_11\,
            carryout => \display2.prescaler_2_cry_12\,
            clk => \N__14237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_13_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13253\,
            in2 => \_gnd_net_\,
            in3 => \N__12897\,
            lcout => \display2.prescalerZ0Z_13\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_12\,
            carryout => \display2.prescaler_2_cry_13\,
            clk => \N__14237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_14_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13155\,
            in2 => \_gnd_net_\,
            in3 => \N__12894\,
            lcout => \display2.prescaler_2_14\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_13\,
            carryout => \display2.prescaler_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNO_0_15_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13952\,
            in2 => \_gnd_net_\,
            in3 => \N__12891\,
            lcout => \display2.prescaler_2_15\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_14\,
            carryout => \display2.prescaler_2_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_16_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13131\,
            in2 => \_gnd_net_\,
            in3 => \N__12888\,
            lcout => \display2.prescalerZ0Z_16\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_15\,
            carryout => \display2.prescaler_2_cry_16\,
            clk => \N__14237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_17_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13143\,
            in2 => \_gnd_net_\,
            in3 => \N__12885\,
            lcout => \display2.prescalerZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \display2.prescaler_2_cry_17\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_18_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13118\,
            in2 => \_gnd_net_\,
            in3 => \N__12882\,
            lcout => \display2.prescalerZ0Z_18\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_17\,
            carryout => \display2.prescaler_2_cry_18\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_19_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12969\,
            in3 => \N__13032\,
            lcout => \display2.prescalerZ0Z_19\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_18\,
            carryout => \display2.prescaler_2_cry_19\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_20_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12993\,
            in2 => \_gnd_net_\,
            in3 => \N__13029\,
            lcout => \display2.prescalerZ0Z_20\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_19\,
            carryout => \display2.prescaler_2_cry_20\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_21_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13002\,
            in2 => \_gnd_net_\,
            in3 => \N__13026\,
            lcout => \display2.prescalerZ0Z_21\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_20\,
            carryout => \display2.prescaler_2_cry_21\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_22_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12984\,
            in3 => \N__13023\,
            lcout => \display2.prescalerZ0Z_22\,
            ltout => OPEN,
            carryin => \display2.prescaler_2_cry_21\,
            carryout => \display2.prescaler_2_cry_22\,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_23_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13016\,
            in2 => \_gnd_net_\,
            in3 => \N__13020\,
            lcout => \display2.prescalerZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNIF8K21_19_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13001\,
            in1 => \N__12992\,
            in2 => \N__12983\,
            in3 => \N__12965\,
            lcout => \display2.prescaler8_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNIDHIG_2_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12956\,
            in1 => \N__12944\,
            in2 => \N__12933\,
            in3 => \N__12917\,
            lcout => \display2.prescaler8_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.digit_posn_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__14032\,
            in2 => \N__13410\,
            in3 => \N__13994\,
            lcout => \display2.digit_posnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_0_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__13995\,
            in1 => \N__13069\,
            in2 => \N__14042\,
            in3 => \N__13103\,
            lcout => \display2.prescalerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_1_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13205\,
            lcout => \display2.prescalerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNI6SG21_10_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13284\,
            in1 => \N__13268\,
            in2 => \N__13257\,
            in3 => \N__13238\,
            lcout => OPEN,
            ltout => \display2.prescaler8_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNI7PO13_1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13227\,
            in1 => \N__13185\,
            in2 => \N__13218\,
            in3 => \N__13215\,
            lcout => \display2.prescaler8_21\,
            ltout => \display2.prescaler8_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNIQNE25_16_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__13990\,
            in1 => \_gnd_net_\,
            in2 => \N__13209\,
            in3 => \N__13057\,
            lcout => \display2.prescaler8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNIHUHP_1_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13154\,
            in1 => \N__13172\,
            in2 => \N__13953\,
            in3 => \N__13204\,
            lcout => \display2.prescaler8_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_9_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__13993\,
            in1 => \N__14031\,
            in2 => \N__13081\,
            in3 => \N__13179\,
            lcout => \display2.prescalerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_14_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__14030\,
            in1 => \N__13991\,
            in2 => \N__13073\,
            in3 => \N__13161\,
            lcout => \display2.prescalerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_RNI4M1U_16_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13142\,
            in1 => \N__13130\,
            in2 => \N__13119\,
            in3 => \N__13102\,
            lcout => \display2.prescaler8_17\,
            ltout => \display2.prescaler8_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.prescaler_15_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__14049\,
            in1 => \N__14036\,
            in2 => \N__13998\,
            in3 => \N__13992\,
            lcout => \display2.prescalerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_0_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \d1.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.digit_data_3_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__13344\,
            in1 => \N__13401\,
            in2 => \N__14465\,
            in3 => \N__13896\,
            lcout => \display2.digit_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.digit_data_2_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__13400\,
            in1 => \N__13343\,
            in2 => \N__14521\,
            in3 => \N__13794\,
            lcout => \display2.digit_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.digit_data_1_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__13346\,
            in1 => \N__13412\,
            in2 => \N__14388\,
            in3 => \N__13683\,
            lcout => \display2.digit_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.digit_data_0_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__13411\,
            in1 => \N__13345\,
            in2 => \N__14331\,
            in3 => \N__13554\,
            lcout => \display2.digit_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.DIGIT_e_0_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13416\,
            lcout => \DIGIT_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14257\,
            ce => \N__13353\,
            sr => \_gnd_net_\
        );

    \d4.sync_0_LC_19_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13323\,
            lcout => \d4.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_0_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000110110"
        )
    port map (
            in0 => \N__14522\,
            in1 => \N__14476\,
            in2 => \N__14423\,
            in3 => \N__14350\,
            lcout => \SEG2_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_5_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100010111"
        )
    port map (
            in0 => \N__14541\,
            in1 => \N__14478\,
            in2 => \N__14405\,
            in3 => \N__14332\,
            lcout => \SEG2_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_2_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__14352\,
            in1 => \N__14524\,
            in2 => \N__14477\,
            in3 => \N__14422\,
            lcout => \SEG2_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_1_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000100111"
        )
    port map (
            in0 => \N__14523\,
            in1 => \N__14461\,
            in2 => \N__14424\,
            in3 => \N__14351\,
            lcout => \SEG2_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_4_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100111011"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__14395\,
            in2 => \N__14484\,
            in3 => \N__14543\,
            lcout => \SEG2_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_3_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000110101"
        )
    port map (
            in0 => \N__14542\,
            in1 => \N__14479\,
            in2 => \N__14406\,
            in3 => \N__14333\,
            lcout => \SEG2_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display2.decoder.SEG_6_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011000110101"
        )
    port map (
            in0 => \N__14544\,
            in1 => \N__14480\,
            in2 => \N__14407\,
            in3 => \N__14335\,
            lcout => \SEG2_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14275\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
