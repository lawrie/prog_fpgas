// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Dec 23 2017 18:12:09

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "servo_tester" view "INTERFACE"

module servo_tester (
    switch_up,
    switch_dn,
    CONTROL_PIN,
    CLK);

    input switch_up;
    input switch_dn;
    output CONTROL_PIN;
    input CLK;

    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4954;
    wire N__4951;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4939;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4924;
    wire N__4921;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4906;
    wire N__4903;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4803;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4793;
    wire N__4792;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4705;
    wire N__4702;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4690;
    wire N__4687;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4675;
    wire N__4672;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4642;
    wire N__4639;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4627;
    wire N__4624;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4591;
    wire N__4590;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4578;
    wire N__4573;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4543;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4507;
    wire N__4506;
    wire N__4505;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4488;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4460;
    wire N__4459;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4441;
    wire N__4440;
    wire N__4439;
    wire N__4434;
    wire N__4431;
    wire N__4430;
    wire N__4429;
    wire N__4428;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4396;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4378;
    wire N__4375;
    wire N__4374;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4354;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4327;
    wire N__4324;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4312;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4294;
    wire N__4291;
    wire N__4290;
    wire N__4289;
    wire N__4286;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4255;
    wire N__4252;
    wire N__4251;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4237;
    wire N__4234;
    wire N__4233;
    wire N__4230;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4207;
    wire N__4204;
    wire N__4203;
    wire N__4202;
    wire N__4199;
    wire N__4194;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4117;
    wire N__4116;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4101;
    wire N__4100;
    wire N__4097;
    wire N__4092;
    wire N__4085;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4074;
    wire N__4073;
    wire N__4070;
    wire N__4063;
    wire N__4060;
    wire N__4053;
    wire N__4050;
    wire N__4043;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4008;
    wire N__4005;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3988;
    wire N__3985;
    wire N__3984;
    wire N__3983;
    wire N__3980;
    wire N__3979;
    wire N__3978;
    wire N__3973;
    wire N__3970;
    wire N__3965;
    wire N__3958;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3922;
    wire N__3921;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3901;
    wire N__3900;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3877;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3856;
    wire N__3855;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3814;
    wire N__3813;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3790;
    wire N__3789;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3769;
    wire N__3768;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3748;
    wire N__3747;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3727;
    wire N__3726;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3703;
    wire N__3702;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3665;
    wire N__3664;
    wire N__3663;
    wire N__3658;
    wire N__3655;
    wire N__3650;
    wire N__3643;
    wire N__3642;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3622;
    wire N__3621;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3517;
    wire N__3514;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3465;
    wire N__3464;
    wire N__3463;
    wire N__3462;
    wire N__3461;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3457;
    wire N__3456;
    wire N__3455;
    wire N__3448;
    wire N__3441;
    wire N__3438;
    wire N__3431;
    wire N__3426;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3399;
    wire N__3398;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3384;
    wire N__3383;
    wire N__3378;
    wire N__3375;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3336;
    wire N__3335;
    wire N__3332;
    wire N__3331;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3315;
    wire N__3310;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2802;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2787;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2771;
    wire N__2766;
    wire N__2761;
    wire N__2760;
    wire N__2759;
    wire N__2758;
    wire N__2755;
    wire N__2748;
    wire N__2743;
    wire N__2740;
    wire N__2739;
    wire N__2738;
    wire N__2735;
    wire N__2730;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2698;
    wire N__2695;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2683;
    wire N__2680;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2665;
    wire N__2662;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire N__2652;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2563;
    wire N__2560;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2548;
    wire N__2545;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2533;
    wire N__2530;
    wire N__2529;
    wire N__2526;
    wire N__2523;
    wire N__2518;
    wire N__2515;
    wire N__2514;
    wire N__2511;
    wire N__2508;
    wire N__2503;
    wire N__2500;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2488;
    wire N__2485;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2475;
    wire N__2470;
    wire N__2467;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2455;
    wire N__2452;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2440;
    wire N__2437;
    wire N__2436;
    wire N__2433;
    wire N__2430;
    wire N__2425;
    wire N__2422;
    wire N__2419;
    wire N__2416;
    wire N__2415;
    wire N__2412;
    wire N__2409;
    wire N__2404;
    wire N__2401;
    wire N__2400;
    wire N__2397;
    wire N__2394;
    wire N__2389;
    wire N__2386;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2374;
    wire N__2371;
    wire N__2370;
    wire N__2367;
    wire N__2364;
    wire N__2359;
    wire N__2356;
    wire N__2355;
    wire N__2352;
    wire N__2349;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2320;
    wire N__2317;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2301;
    wire N__2300;
    wire N__2297;
    wire N__2292;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_11_0_;
    wire \p.prescaler12_0 ;
    wire \p.prescaler12_1 ;
    wire \p.prescaler12_2 ;
    wire \p.prescaler12_3 ;
    wire \p.prescaler12_4 ;
    wire \p.prescaler12_5 ;
    wire \p.prescaler12 ;
    wire \p.prescaler12_THRU_CO ;
    wire \p.prescaler12_4_and ;
    wire \p.prescaler12_2_and ;
    wire \p.prescaler12_6_and ;
    wire \p.prescaler12_5_and ;
    wire \p.prescaler12_3_and ;
    wire \p.prescaler12_1_and ;
    wire bfn_2_11_0_;
    wire \p.prescalerZ0Z_2 ;
    wire \p.prescaler_1_cry_1_THRU_CO ;
    wire \p.prescaler_1_cry_1 ;
    wire \p.prescalerZ0Z_3 ;
    wire \p.prescaler_1_cry_2 ;
    wire \p.prescalerZ0Z_4 ;
    wire \p.prescaler_1_cry_3 ;
    wire \p.prescaler_1_cry_4 ;
    wire \p.prescaler_1_cry_5 ;
    wire \p.prescalerZ0Z_7 ;
    wire \p.prescaler_1_cry_6 ;
    wire \p.prescalerZ0Z_8 ;
    wire \p.prescaler_1_cry_7 ;
    wire \p.prescaler_1_cry_8 ;
    wire \p.prescalerZ0Z_9 ;
    wire bfn_2_12_0_;
    wire \p.prescalerZ0Z_10 ;
    wire \p.prescaler_1_cry_9 ;
    wire \p.prescalerZ0Z_11 ;
    wire \p.prescaler_1_cry_10 ;
    wire \p.prescalerZ0Z_12 ;
    wire \p.prescaler_1_cry_11 ;
    wire \p.prescalerZ0Z_13 ;
    wire \p.prescaler_1_cry_12 ;
    wire \p.prescalerZ0Z_14 ;
    wire \p.prescaler_1_cry_13 ;
    wire \p.prescalerZ0Z_15 ;
    wire \p.prescaler_1_cry_14 ;
    wire \p.prescalerZ0Z_16 ;
    wire \p.prescaler_1_cry_15 ;
    wire \p.prescaler_1_cry_16 ;
    wire \p.prescalerZ0Z_17 ;
    wire bfn_2_13_0_;
    wire \p.prescalerZ0Z_18 ;
    wire \p.prescaler_1_cry_17 ;
    wire \p.prescalerZ0Z_19 ;
    wire \p.prescaler_1_cry_18 ;
    wire \p.prescalerZ0Z_20 ;
    wire \p.prescaler_1_cry_19 ;
    wire \p.prescalerZ0Z_21 ;
    wire \p.prescaler_1_cry_20 ;
    wire \p.prescalerZ0Z_22 ;
    wire \p.prescaler_1_cry_21 ;
    wire \p.prescalerZ0Z_23 ;
    wire \p.prescaler_1_cry_22 ;
    wire \p.prescalerZ0Z_24 ;
    wire \p.prescaler_1_cry_23 ;
    wire \p.prescaler_1_cry_24 ;
    wire \p.prescalerZ0Z_25 ;
    wire bfn_2_14_0_;
    wire \p.prescaler_1_cry_25 ;
    wire \p.prescalerZ0Z_26 ;
    wire \p.prescaler12_0_and ;
    wire \p.prescaler_1_cry_5_THRU_CO ;
    wire \p.prescalerZ0Z_6 ;
    wire \p.prescaler_1_cry_4_THRU_CO ;
    wire \p.prescalerZ0Z_5 ;
    wire \p.prescalerZ0Z_0 ;
    wire \p.prescalerZ0Z_1 ;
    wire bfn_7_8_0_;
    wire state_RNIPC4P3;
    wire un1_pulse_len_cry_2;
    wire un1_pulse_len_cry_3;
    wire un1_pulse_len_cry_4;
    wire un1_pulse_len_cry_5;
    wire un1_pulse_len_cry_6;
    wire state_RNIPC4P3_6;
    wire un1_pulse_len_cry_7;
    wire un1_pulse_len_cry_8;
    wire un1_pulse_len_cry_9;
    wire bfn_7_9_0_;
    wire un1_pulse_len_cry_10;
    wire un1_pulse_len_cry_11;
    wire un1_pulse_len_cry_12;
    wire un1_pulse_len_cry_13;
    wire un1_pulse_len_cry_14;
    wire state_RNIPC4P3_4;
    wire state_RNIPC4P3_7;
    wire \p.count_i_2 ;
    wire bfn_7_10_0_;
    wire pulse_lenZ0Z_3;
    wire \p.count_i_3 ;
    wire \p.CONTROL_PIN_2_cry_2 ;
    wire pulse_lenZ0Z_4;
    wire \p.count_i_4 ;
    wire \p.CONTROL_PIN_2_cry_3 ;
    wire pulse_lenZ0Z_5;
    wire \p.count_i_5 ;
    wire \p.CONTROL_PIN_2_cry_4 ;
    wire pulse_lenZ0Z_6;
    wire \p.count_i_6 ;
    wire \p.CONTROL_PIN_2_cry_5 ;
    wire pulse_lenZ0Z_7;
    wire \p.count_i_7 ;
    wire \p.CONTROL_PIN_2_cry_6 ;
    wire pulse_lenZ0Z_8;
    wire \p.count_i_8 ;
    wire \p.CONTROL_PIN_2_cry_7 ;
    wire pulse_lenZ0Z_9;
    wire \p.count_i_9 ;
    wire \p.CONTROL_PIN_2_cry_8 ;
    wire \p.CONTROL_PIN_2_cry_9 ;
    wire pulse_lenZ0Z_10;
    wire \p.count_i_10 ;
    wire bfn_7_11_0_;
    wire pulse_lenZ0Z_11;
    wire \p.count_i_11 ;
    wire \p.CONTROL_PIN_2_cry_10 ;
    wire pulse_lenZ0Z_12;
    wire \p.count_i_12 ;
    wire \p.CONTROL_PIN_2_cry_11 ;
    wire pulse_lenZ0Z_13;
    wire \p.count_i_13 ;
    wire \p.CONTROL_PIN_2_cry_12 ;
    wire pulse_lenZ0Z_14;
    wire \p.count_i_14 ;
    wire \p.CONTROL_PIN_2_cry_13 ;
    wire pulse_lenZ0Z_15;
    wire \p.count_i_15 ;
    wire \p.CONTROL_PIN_2_cry_14 ;
    wire \p.CONTROL_PIN_2 ;
    wire CONTROL_PIN_c;
    wire bfn_7_12_0_;
    wire \p.count_1_cry_1 ;
    wire \p.count_1_cry_2 ;
    wire \p.count_1_cry_3 ;
    wire \p.count_1_cry_4 ;
    wire \p.count_1_cry_5 ;
    wire \p.count_1_cry_6 ;
    wire \p.count_1_cry_7 ;
    wire \p.count_1_cry_8 ;
    wire bfn_7_13_0_;
    wire \p.count_1_cry_9 ;
    wire \p.count_1_cry_10 ;
    wire \p.count_1_cry_11 ;
    wire \p.count_1_cry_12 ;
    wire \p.count_1_cry_13 ;
    wire \p.count_1_cry_14 ;
    wire state_RNIPC4P3_0;
    wire state_RNIPC4P3_2;
    wire \d2.trans_up_1_12_cascade_ ;
    wire \d2.trans_up_1_sx_cascade_ ;
    wire d2_trans_up_1_cascade_;
    wire pulse_lenZ0Z_2;
    wire s_dn_i_cascade_;
    wire un1_pulse_len_cry_2_c_RNOZ0;
    wire state_RNIPC4P3_3;
    wire state_RNIU5D07;
    wire state_RNIPC4P3_1;
    wire state_RNIPC4P3_8;
    wire d2_trans_up_1;
    wire state_RNIPC4P3_5;
    wire \d1.count_RNI2PCEZ0Z_3_cascade_ ;
    wire \d1.trans_up_1_14_cascade_ ;
    wire s_up;
    wire s_up_cascade_;
    wire s_dn_i;
    wire state_RNIU5D07_0;
    wire \d1.trans_up_1_11 ;
    wire \d1.trans_up_1_13_sx_cascade_ ;
    wire \d1.trans_up_1_14 ;
    wire \d1.trans_up_1_13_cascade_ ;
    wire \d1.trans_up_1_12 ;
    wire \d1.trans_up_1_9 ;
    wire \d1.trans_up_sx ;
    wire \d1.stateZ0 ;
    wire \d1.syncZ0Z_1 ;
    wire \d1.idle_i ;
    wire \p.countZ0Z_14 ;
    wire \p.countZ0Z_8 ;
    wire \p.countZ0Z_15 ;
    wire \p.countZ0Z_6 ;
    wire \p.countZ0Z_12 ;
    wire \p.countZ0Z_7 ;
    wire \p.countZ0Z_13 ;
    wire \p.countZ0Z_5 ;
    wire \p.countZ0Z_10 ;
    wire \p.countZ0Z_9 ;
    wire \p.countZ0Z_11 ;
    wire \p.countZ0Z_4 ;
    wire \p.count10_11 ;
    wire \p.count10_10 ;
    wire \p.count10_8_cascade_ ;
    wire \p.count10 ;
    wire \p.countZ0Z_3 ;
    wire \p.countZ0Z_2 ;
    wire \p.count10_9 ;
    wire \d2.trans_up_1_11 ;
    wire \d2.trans_up_1_10 ;
    wire \d2.trans_up_1_9 ;
    wire \d2.count_RNI237Z0Z_11 ;
    wire switch_dn_c;
    wire \d2.syncZ0Z_0 ;
    wire \d2.syncZ0Z_1 ;
    wire d2_state;
    wire \d2.idle_i ;
    wire \d1.countZ0Z_1 ;
    wire \d1.countZ0Z_0 ;
    wire bfn_9_9_0_;
    wire \d1.countZ0Z_2 ;
    wire \d1.un3_count_cry_1 ;
    wire \d1.countZ0Z_3 ;
    wire \d1.un3_count_cry_2 ;
    wire \d1.countZ0Z_4 ;
    wire \d1.un3_count_cry_3 ;
    wire \d1.countZ0Z_5 ;
    wire \d1.un3_count_cry_4 ;
    wire \d1.countZ0Z_6 ;
    wire \d1.un3_count_cry_5 ;
    wire \d1.countZ0Z_7 ;
    wire \d1.un3_count_cry_6 ;
    wire \d1.countZ0Z_8 ;
    wire \d1.un3_count_cry_7 ;
    wire \d1.un3_count_cry_8 ;
    wire \d1.countZ0Z_9 ;
    wire bfn_9_10_0_;
    wire \d1.countZ0Z_10 ;
    wire \d1.un3_count_cry_9 ;
    wire \d1.countZ0Z_11 ;
    wire \d1.un3_count_cry_10 ;
    wire \d1.countZ0Z_12 ;
    wire \d1.un3_count_cry_11 ;
    wire \d1.countZ0Z_13 ;
    wire \d1.un3_count_cry_12 ;
    wire \d1.countZ0Z_14 ;
    wire \d1.un3_count_cry_13 ;
    wire \d1.countZ0Z_15 ;
    wire \d1.un3_count_cry_14 ;
    wire \d1.un3_count_cry_15 ;
    wire \d1.countZ0Z_16 ;
    wire \d1.idle_i_g ;
    wire \p.countZ0Z_1 ;
    wire \p.countZ0Z_0 ;
    wire \p.prescaler12_g ;
    wire \d2.countZ0Z_0 ;
    wire \d2.countZ0Z_1 ;
    wire bfn_9_14_0_;
    wire \d2.countZ0Z_2 ;
    wire \d2.un3_count_cry_1 ;
    wire \d2.countZ0Z_3 ;
    wire \d2.un3_count_cry_2 ;
    wire \d2.countZ0Z_4 ;
    wire \d2.un3_count_cry_3 ;
    wire \d2.countZ0Z_5 ;
    wire \d2.un3_count_cry_4 ;
    wire \d2.countZ0Z_6 ;
    wire \d2.un3_count_cry_5 ;
    wire \d2.countZ0Z_7 ;
    wire \d2.un3_count_cry_6 ;
    wire \d2.countZ0Z_8 ;
    wire \d2.un3_count_cry_7 ;
    wire \d2.un3_count_cry_8 ;
    wire \d2.countZ0Z_9 ;
    wire bfn_9_15_0_;
    wire \d2.countZ0Z_10 ;
    wire \d2.un3_count_cry_9 ;
    wire \d2.countZ0Z_11 ;
    wire \d2.un3_count_cry_10 ;
    wire \d2.countZ0Z_12 ;
    wire \d2.un3_count_cry_11 ;
    wire \d2.countZ0Z_13 ;
    wire \d2.un3_count_cry_12 ;
    wire \d2.countZ0Z_14 ;
    wire \d2.un3_count_cry_13 ;
    wire \d2.countZ0Z_15 ;
    wire \d2.un3_count_cry_14 ;
    wire \d2.un3_count_cry_15 ;
    wire \d2.countZ0Z_16 ;
    wire \d2.idle_i_g ;
    wire switch_up_c;
    wire \d1.syncZ0Z_0 ;
    wire CLK_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5000),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__5002),
            .DIN(N__5001),
            .DOUT(N__5000),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__5002),
            .PADOUT(N__5001),
            .PADIN(N__5000),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD CONTROL_PIN_obuf_iopad (
            .OE(N__4991),
            .DIN(N__4990),
            .DOUT(N__4989),
            .PACKAGEPIN(CONTROL_PIN));
    defparam CONTROL_PIN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONTROL_PIN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONTROL_PIN_obuf_preio (
            .PADOEN(N__4991),
            .PADOUT(N__4990),
            .PADIN(N__4989),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3235),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_dn_ibuf_iopad (
            .OE(N__4982),
            .DIN(N__4981),
            .DOUT(N__4980),
            .PACKAGEPIN(switch_dn));
    defparam switch_dn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_dn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_dn_ibuf_preio (
            .PADOEN(N__4982),
            .PADOUT(N__4981),
            .PADIN(N__4980),
            .CLOCKENABLE(),
            .DIN0(switch_dn_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_up_ibuf_iopad (
            .OE(N__4973),
            .DIN(N__4972),
            .DOUT(N__4971),
            .PACKAGEPIN(switch_up));
    defparam switch_up_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_up_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_up_ibuf_preio (
            .PADOEN(N__4973),
            .PADOUT(N__4972),
            .PADIN(N__4971),
            .CLOCKENABLE(),
            .DIN0(switch_up_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1092 (
            .O(N__4954),
            .I(\d2.un3_count_cry_9 ));
    InMux I__1091 (
            .O(N__4951),
            .I(N__4947));
    InMux I__1090 (
            .O(N__4950),
            .I(N__4944));
    LocalMux I__1089 (
            .O(N__4947),
            .I(\d2.countZ0Z_11 ));
    LocalMux I__1088 (
            .O(N__4944),
            .I(\d2.countZ0Z_11 ));
    InMux I__1087 (
            .O(N__4939),
            .I(\d2.un3_count_cry_10 ));
    InMux I__1086 (
            .O(N__4936),
            .I(N__4932));
    InMux I__1085 (
            .O(N__4935),
            .I(N__4929));
    LocalMux I__1084 (
            .O(N__4932),
            .I(\d2.countZ0Z_12 ));
    LocalMux I__1083 (
            .O(N__4929),
            .I(\d2.countZ0Z_12 ));
    InMux I__1082 (
            .O(N__4924),
            .I(\d2.un3_count_cry_11 ));
    CascadeMux I__1081 (
            .O(N__4921),
            .I(N__4917));
    InMux I__1080 (
            .O(N__4920),
            .I(N__4914));
    InMux I__1079 (
            .O(N__4917),
            .I(N__4911));
    LocalMux I__1078 (
            .O(N__4914),
            .I(\d2.countZ0Z_13 ));
    LocalMux I__1077 (
            .O(N__4911),
            .I(\d2.countZ0Z_13 ));
    InMux I__1076 (
            .O(N__4906),
            .I(\d2.un3_count_cry_12 ));
    InMux I__1075 (
            .O(N__4903),
            .I(N__4899));
    InMux I__1074 (
            .O(N__4902),
            .I(N__4896));
    LocalMux I__1073 (
            .O(N__4899),
            .I(\d2.countZ0Z_14 ));
    LocalMux I__1072 (
            .O(N__4896),
            .I(\d2.countZ0Z_14 ));
    InMux I__1071 (
            .O(N__4891),
            .I(\d2.un3_count_cry_13 ));
    InMux I__1070 (
            .O(N__4888),
            .I(N__4884));
    InMux I__1069 (
            .O(N__4887),
            .I(N__4881));
    LocalMux I__1068 (
            .O(N__4884),
            .I(\d2.countZ0Z_15 ));
    LocalMux I__1067 (
            .O(N__4881),
            .I(\d2.countZ0Z_15 ));
    InMux I__1066 (
            .O(N__4876),
            .I(\d2.un3_count_cry_14 ));
    InMux I__1065 (
            .O(N__4873),
            .I(\d2.un3_count_cry_15 ));
    InMux I__1064 (
            .O(N__4870),
            .I(N__4866));
    InMux I__1063 (
            .O(N__4869),
            .I(N__4863));
    LocalMux I__1062 (
            .O(N__4866),
            .I(N__4860));
    LocalMux I__1061 (
            .O(N__4863),
            .I(\d2.countZ0Z_16 ));
    Odrv4 I__1060 (
            .O(N__4860),
            .I(\d2.countZ0Z_16 ));
    SRMux I__1059 (
            .O(N__4855),
            .I(N__4846));
    SRMux I__1058 (
            .O(N__4854),
            .I(N__4846));
    SRMux I__1057 (
            .O(N__4853),
            .I(N__4846));
    GlobalMux I__1056 (
            .O(N__4846),
            .I(N__4843));
    gio2CtrlBuf I__1055 (
            .O(N__4843),
            .I(\d2.idle_i_g ));
    InMux I__1054 (
            .O(N__4840),
            .I(N__4837));
    LocalMux I__1053 (
            .O(N__4837),
            .I(N__4834));
    Span12Mux_h I__1052 (
            .O(N__4834),
            .I(N__4831));
    Span12Mux_v I__1051 (
            .O(N__4831),
            .I(N__4828));
    Span12Mux_h I__1050 (
            .O(N__4828),
            .I(N__4825));
    Odrv12 I__1049 (
            .O(N__4825),
            .I(switch_up_c));
    InMux I__1048 (
            .O(N__4822),
            .I(N__4819));
    LocalMux I__1047 (
            .O(N__4819),
            .I(N__4816));
    Odrv12 I__1046 (
            .O(N__4816),
            .I(\d1.syncZ0Z_0 ));
    ClkMux I__1045 (
            .O(N__4813),
            .I(N__4738));
    ClkMux I__1044 (
            .O(N__4812),
            .I(N__4738));
    ClkMux I__1043 (
            .O(N__4811),
            .I(N__4738));
    ClkMux I__1042 (
            .O(N__4810),
            .I(N__4738));
    ClkMux I__1041 (
            .O(N__4809),
            .I(N__4738));
    ClkMux I__1040 (
            .O(N__4808),
            .I(N__4738));
    ClkMux I__1039 (
            .O(N__4807),
            .I(N__4738));
    ClkMux I__1038 (
            .O(N__4806),
            .I(N__4738));
    ClkMux I__1037 (
            .O(N__4805),
            .I(N__4738));
    ClkMux I__1036 (
            .O(N__4804),
            .I(N__4738));
    ClkMux I__1035 (
            .O(N__4803),
            .I(N__4738));
    ClkMux I__1034 (
            .O(N__4802),
            .I(N__4738));
    ClkMux I__1033 (
            .O(N__4801),
            .I(N__4738));
    ClkMux I__1032 (
            .O(N__4800),
            .I(N__4738));
    ClkMux I__1031 (
            .O(N__4799),
            .I(N__4738));
    ClkMux I__1030 (
            .O(N__4798),
            .I(N__4738));
    ClkMux I__1029 (
            .O(N__4797),
            .I(N__4738));
    ClkMux I__1028 (
            .O(N__4796),
            .I(N__4738));
    ClkMux I__1027 (
            .O(N__4795),
            .I(N__4738));
    ClkMux I__1026 (
            .O(N__4794),
            .I(N__4738));
    ClkMux I__1025 (
            .O(N__4793),
            .I(N__4738));
    ClkMux I__1024 (
            .O(N__4792),
            .I(N__4738));
    ClkMux I__1023 (
            .O(N__4791),
            .I(N__4738));
    ClkMux I__1022 (
            .O(N__4790),
            .I(N__4738));
    ClkMux I__1021 (
            .O(N__4789),
            .I(N__4738));
    GlobalMux I__1020 (
            .O(N__4738),
            .I(N__4735));
    gio2CtrlBuf I__1019 (
            .O(N__4735),
            .I(CLK_c_g));
    InMux I__1018 (
            .O(N__4732),
            .I(N__4728));
    InMux I__1017 (
            .O(N__4731),
            .I(N__4725));
    LocalMux I__1016 (
            .O(N__4728),
            .I(\d2.countZ0Z_2 ));
    LocalMux I__1015 (
            .O(N__4725),
            .I(\d2.countZ0Z_2 ));
    InMux I__1014 (
            .O(N__4720),
            .I(\d2.un3_count_cry_1 ));
    InMux I__1013 (
            .O(N__4717),
            .I(N__4713));
    InMux I__1012 (
            .O(N__4716),
            .I(N__4710));
    LocalMux I__1011 (
            .O(N__4713),
            .I(\d2.countZ0Z_3 ));
    LocalMux I__1010 (
            .O(N__4710),
            .I(\d2.countZ0Z_3 ));
    InMux I__1009 (
            .O(N__4705),
            .I(\d2.un3_count_cry_2 ));
    InMux I__1008 (
            .O(N__4702),
            .I(N__4698));
    InMux I__1007 (
            .O(N__4701),
            .I(N__4695));
    LocalMux I__1006 (
            .O(N__4698),
            .I(\d2.countZ0Z_4 ));
    LocalMux I__1005 (
            .O(N__4695),
            .I(\d2.countZ0Z_4 ));
    InMux I__1004 (
            .O(N__4690),
            .I(\d2.un3_count_cry_3 ));
    InMux I__1003 (
            .O(N__4687),
            .I(N__4683));
    InMux I__1002 (
            .O(N__4686),
            .I(N__4680));
    LocalMux I__1001 (
            .O(N__4683),
            .I(\d2.countZ0Z_5 ));
    LocalMux I__1000 (
            .O(N__4680),
            .I(\d2.countZ0Z_5 ));
    InMux I__999 (
            .O(N__4675),
            .I(\d2.un3_count_cry_4 ));
    CascadeMux I__998 (
            .O(N__4672),
            .I(N__4668));
    InMux I__997 (
            .O(N__4671),
            .I(N__4665));
    InMux I__996 (
            .O(N__4668),
            .I(N__4662));
    LocalMux I__995 (
            .O(N__4665),
            .I(\d2.countZ0Z_6 ));
    LocalMux I__994 (
            .O(N__4662),
            .I(\d2.countZ0Z_6 ));
    InMux I__993 (
            .O(N__4657),
            .I(\d2.un3_count_cry_5 ));
    InMux I__992 (
            .O(N__4654),
            .I(N__4650));
    InMux I__991 (
            .O(N__4653),
            .I(N__4647));
    LocalMux I__990 (
            .O(N__4650),
            .I(\d2.countZ0Z_7 ));
    LocalMux I__989 (
            .O(N__4647),
            .I(\d2.countZ0Z_7 ));
    InMux I__988 (
            .O(N__4642),
            .I(\d2.un3_count_cry_6 ));
    InMux I__987 (
            .O(N__4639),
            .I(N__4635));
    InMux I__986 (
            .O(N__4638),
            .I(N__4632));
    LocalMux I__985 (
            .O(N__4635),
            .I(\d2.countZ0Z_8 ));
    LocalMux I__984 (
            .O(N__4632),
            .I(\d2.countZ0Z_8 ));
    InMux I__983 (
            .O(N__4627),
            .I(\d2.un3_count_cry_7 ));
    InMux I__982 (
            .O(N__4624),
            .I(N__4620));
    InMux I__981 (
            .O(N__4623),
            .I(N__4617));
    LocalMux I__980 (
            .O(N__4620),
            .I(\d2.countZ0Z_9 ));
    LocalMux I__979 (
            .O(N__4617),
            .I(\d2.countZ0Z_9 ));
    InMux I__978 (
            .O(N__4612),
            .I(bfn_9_15_0_));
    CascadeMux I__977 (
            .O(N__4609),
            .I(N__4606));
    InMux I__976 (
            .O(N__4606),
            .I(N__4602));
    InMux I__975 (
            .O(N__4605),
            .I(N__4599));
    LocalMux I__974 (
            .O(N__4602),
            .I(N__4596));
    LocalMux I__973 (
            .O(N__4599),
            .I(\d2.countZ0Z_10 ));
    Odrv4 I__972 (
            .O(N__4596),
            .I(\d2.countZ0Z_10 ));
    CascadeMux I__971 (
            .O(N__4591),
            .I(N__4586));
    InMux I__970 (
            .O(N__4590),
            .I(N__4583));
    InMux I__969 (
            .O(N__4589),
            .I(N__4578));
    InMux I__968 (
            .O(N__4586),
            .I(N__4578));
    LocalMux I__967 (
            .O(N__4583),
            .I(\d1.countZ0Z_12 ));
    LocalMux I__966 (
            .O(N__4578),
            .I(\d1.countZ0Z_12 ));
    InMux I__965 (
            .O(N__4573),
            .I(\d1.un3_count_cry_11 ));
    InMux I__964 (
            .O(N__4570),
            .I(N__4566));
    InMux I__963 (
            .O(N__4569),
            .I(N__4563));
    LocalMux I__962 (
            .O(N__4566),
            .I(\d1.countZ0Z_13 ));
    LocalMux I__961 (
            .O(N__4563),
            .I(\d1.countZ0Z_13 ));
    InMux I__960 (
            .O(N__4558),
            .I(\d1.un3_count_cry_12 ));
    InMux I__959 (
            .O(N__4555),
            .I(N__4551));
    InMux I__958 (
            .O(N__4554),
            .I(N__4548));
    LocalMux I__957 (
            .O(N__4551),
            .I(\d1.countZ0Z_14 ));
    LocalMux I__956 (
            .O(N__4548),
            .I(\d1.countZ0Z_14 ));
    InMux I__955 (
            .O(N__4543),
            .I(\d1.un3_count_cry_13 ));
    InMux I__954 (
            .O(N__4540),
            .I(N__4536));
    InMux I__953 (
            .O(N__4539),
            .I(N__4533));
    LocalMux I__952 (
            .O(N__4536),
            .I(\d1.countZ0Z_15 ));
    LocalMux I__951 (
            .O(N__4533),
            .I(\d1.countZ0Z_15 ));
    InMux I__950 (
            .O(N__4528),
            .I(\d1.un3_count_cry_14 ));
    InMux I__949 (
            .O(N__4525),
            .I(\d1.un3_count_cry_15 ));
    CascadeMux I__948 (
            .O(N__4522),
            .I(N__4518));
    InMux I__947 (
            .O(N__4521),
            .I(N__4515));
    InMux I__946 (
            .O(N__4518),
            .I(N__4512));
    LocalMux I__945 (
            .O(N__4515),
            .I(\d1.countZ0Z_16 ));
    LocalMux I__944 (
            .O(N__4512),
            .I(\d1.countZ0Z_16 ));
    SRMux I__943 (
            .O(N__4507),
            .I(N__4498));
    SRMux I__942 (
            .O(N__4506),
            .I(N__4498));
    SRMux I__941 (
            .O(N__4505),
            .I(N__4498));
    GlobalMux I__940 (
            .O(N__4498),
            .I(N__4495));
    gio2CtrlBuf I__939 (
            .O(N__4495),
            .I(\d1.idle_i_g ));
    CascadeMux I__938 (
            .O(N__4492),
            .I(N__4489));
    InMux I__937 (
            .O(N__4489),
            .I(N__4484));
    CascadeMux I__936 (
            .O(N__4488),
            .I(N__4481));
    InMux I__935 (
            .O(N__4487),
            .I(N__4478));
    LocalMux I__934 (
            .O(N__4484),
            .I(N__4475));
    InMux I__933 (
            .O(N__4481),
            .I(N__4472));
    LocalMux I__932 (
            .O(N__4478),
            .I(\p.countZ0Z_1 ));
    Odrv4 I__931 (
            .O(N__4475),
            .I(\p.countZ0Z_1 ));
    LocalMux I__930 (
            .O(N__4472),
            .I(\p.countZ0Z_1 ));
    InMux I__929 (
            .O(N__4465),
            .I(N__4460));
    InMux I__928 (
            .O(N__4464),
            .I(N__4454));
    InMux I__927 (
            .O(N__4463),
            .I(N__4454));
    LocalMux I__926 (
            .O(N__4460),
            .I(N__4451));
    InMux I__925 (
            .O(N__4459),
            .I(N__4448));
    LocalMux I__924 (
            .O(N__4454),
            .I(\p.countZ0Z_0 ));
    Odrv4 I__923 (
            .O(N__4451),
            .I(\p.countZ0Z_0 ));
    LocalMux I__922 (
            .O(N__4448),
            .I(\p.countZ0Z_0 ));
    InMux I__921 (
            .O(N__4441),
            .I(N__4434));
    InMux I__920 (
            .O(N__4440),
            .I(N__4434));
    InMux I__919 (
            .O(N__4439),
            .I(N__4431));
    LocalMux I__918 (
            .O(N__4434),
            .I(N__4424));
    LocalMux I__917 (
            .O(N__4431),
            .I(N__4421));
    CEMux I__916 (
            .O(N__4430),
            .I(N__4408));
    CEMux I__915 (
            .O(N__4429),
            .I(N__4408));
    CEMux I__914 (
            .O(N__4428),
            .I(N__4408));
    CEMux I__913 (
            .O(N__4427),
            .I(N__4408));
    Glb2LocalMux I__912 (
            .O(N__4424),
            .I(N__4408));
    Glb2LocalMux I__911 (
            .O(N__4421),
            .I(N__4408));
    GlobalMux I__910 (
            .O(N__4408),
            .I(N__4405));
    gio2CtrlBuf I__909 (
            .O(N__4405),
            .I(\p.prescaler12_g ));
    InMux I__908 (
            .O(N__4402),
            .I(N__4397));
    InMux I__907 (
            .O(N__4401),
            .I(N__4391));
    InMux I__906 (
            .O(N__4400),
            .I(N__4391));
    LocalMux I__905 (
            .O(N__4397),
            .I(N__4388));
    InMux I__904 (
            .O(N__4396),
            .I(N__4385));
    LocalMux I__903 (
            .O(N__4391),
            .I(\d2.countZ0Z_0 ));
    Odrv12 I__902 (
            .O(N__4388),
            .I(\d2.countZ0Z_0 ));
    LocalMux I__901 (
            .O(N__4385),
            .I(\d2.countZ0Z_0 ));
    CascadeMux I__900 (
            .O(N__4378),
            .I(N__4375));
    InMux I__899 (
            .O(N__4375),
            .I(N__4371));
    InMux I__898 (
            .O(N__4374),
            .I(N__4367));
    LocalMux I__897 (
            .O(N__4371),
            .I(N__4364));
    InMux I__896 (
            .O(N__4370),
            .I(N__4361));
    LocalMux I__895 (
            .O(N__4367),
            .I(\d2.countZ0Z_1 ));
    Odrv12 I__894 (
            .O(N__4364),
            .I(\d2.countZ0Z_1 ));
    LocalMux I__893 (
            .O(N__4361),
            .I(\d2.countZ0Z_1 ));
    InMux I__892 (
            .O(N__4354),
            .I(N__4350));
    InMux I__891 (
            .O(N__4353),
            .I(N__4347));
    LocalMux I__890 (
            .O(N__4350),
            .I(\d1.countZ0Z_3 ));
    LocalMux I__889 (
            .O(N__4347),
            .I(\d1.countZ0Z_3 ));
    InMux I__888 (
            .O(N__4342),
            .I(\d1.un3_count_cry_2 ));
    InMux I__887 (
            .O(N__4339),
            .I(N__4335));
    InMux I__886 (
            .O(N__4338),
            .I(N__4332));
    LocalMux I__885 (
            .O(N__4335),
            .I(\d1.countZ0Z_4 ));
    LocalMux I__884 (
            .O(N__4332),
            .I(\d1.countZ0Z_4 ));
    InMux I__883 (
            .O(N__4327),
            .I(\d1.un3_count_cry_3 ));
    InMux I__882 (
            .O(N__4324),
            .I(N__4320));
    InMux I__881 (
            .O(N__4323),
            .I(N__4317));
    LocalMux I__880 (
            .O(N__4320),
            .I(\d1.countZ0Z_5 ));
    LocalMux I__879 (
            .O(N__4317),
            .I(\d1.countZ0Z_5 ));
    InMux I__878 (
            .O(N__4312),
            .I(\d1.un3_count_cry_4 ));
    CascadeMux I__877 (
            .O(N__4309),
            .I(N__4305));
    InMux I__876 (
            .O(N__4308),
            .I(N__4302));
    InMux I__875 (
            .O(N__4305),
            .I(N__4299));
    LocalMux I__874 (
            .O(N__4302),
            .I(\d1.countZ0Z_6 ));
    LocalMux I__873 (
            .O(N__4299),
            .I(\d1.countZ0Z_6 ));
    InMux I__872 (
            .O(N__4294),
            .I(\d1.un3_count_cry_5 ));
    InMux I__871 (
            .O(N__4291),
            .I(N__4286));
    InMux I__870 (
            .O(N__4290),
            .I(N__4281));
    InMux I__869 (
            .O(N__4289),
            .I(N__4281));
    LocalMux I__868 (
            .O(N__4286),
            .I(\d1.countZ0Z_7 ));
    LocalMux I__867 (
            .O(N__4281),
            .I(\d1.countZ0Z_7 ));
    InMux I__866 (
            .O(N__4276),
            .I(\d1.un3_count_cry_6 ));
    InMux I__865 (
            .O(N__4273),
            .I(N__4268));
    InMux I__864 (
            .O(N__4272),
            .I(N__4265));
    InMux I__863 (
            .O(N__4271),
            .I(N__4262));
    LocalMux I__862 (
            .O(N__4268),
            .I(\d1.countZ0Z_8 ));
    LocalMux I__861 (
            .O(N__4265),
            .I(\d1.countZ0Z_8 ));
    LocalMux I__860 (
            .O(N__4262),
            .I(\d1.countZ0Z_8 ));
    InMux I__859 (
            .O(N__4255),
            .I(\d1.un3_count_cry_7 ));
    InMux I__858 (
            .O(N__4252),
            .I(N__4247));
    InMux I__857 (
            .O(N__4251),
            .I(N__4242));
    InMux I__856 (
            .O(N__4250),
            .I(N__4242));
    LocalMux I__855 (
            .O(N__4247),
            .I(\d1.countZ0Z_9 ));
    LocalMux I__854 (
            .O(N__4242),
            .I(\d1.countZ0Z_9 ));
    InMux I__853 (
            .O(N__4237),
            .I(bfn_9_10_0_));
    CascadeMux I__852 (
            .O(N__4234),
            .I(N__4230));
    CascadeMux I__851 (
            .O(N__4233),
            .I(N__4226));
    InMux I__850 (
            .O(N__4230),
            .I(N__4223));
    InMux I__849 (
            .O(N__4229),
            .I(N__4220));
    InMux I__848 (
            .O(N__4226),
            .I(N__4217));
    LocalMux I__847 (
            .O(N__4223),
            .I(N__4214));
    LocalMux I__846 (
            .O(N__4220),
            .I(\d1.countZ0Z_10 ));
    LocalMux I__845 (
            .O(N__4217),
            .I(\d1.countZ0Z_10 ));
    Odrv4 I__844 (
            .O(N__4214),
            .I(\d1.countZ0Z_10 ));
    InMux I__843 (
            .O(N__4207),
            .I(\d1.un3_count_cry_9 ));
    InMux I__842 (
            .O(N__4204),
            .I(N__4199));
    InMux I__841 (
            .O(N__4203),
            .I(N__4194));
    InMux I__840 (
            .O(N__4202),
            .I(N__4194));
    LocalMux I__839 (
            .O(N__4199),
            .I(\d1.countZ0Z_11 ));
    LocalMux I__838 (
            .O(N__4194),
            .I(\d1.countZ0Z_11 ));
    InMux I__837 (
            .O(N__4189),
            .I(\d1.un3_count_cry_10 ));
    InMux I__836 (
            .O(N__4186),
            .I(N__4183));
    LocalMux I__835 (
            .O(N__4183),
            .I(N__4180));
    Span4Mux_v I__834 (
            .O(N__4180),
            .I(N__4177));
    Odrv4 I__833 (
            .O(N__4177),
            .I(\d2.trans_up_1_9 ));
    InMux I__832 (
            .O(N__4174),
            .I(N__4171));
    LocalMux I__831 (
            .O(N__4171),
            .I(N__4168));
    Span4Mux_v I__830 (
            .O(N__4168),
            .I(N__4165));
    Span4Mux_v I__829 (
            .O(N__4165),
            .I(N__4162));
    Odrv4 I__828 (
            .O(N__4162),
            .I(\d2.count_RNI237Z0Z_11 ));
    InMux I__827 (
            .O(N__4159),
            .I(N__4156));
    LocalMux I__826 (
            .O(N__4156),
            .I(N__4153));
    Span4Mux_v I__825 (
            .O(N__4153),
            .I(N__4150));
    Span4Mux_h I__824 (
            .O(N__4150),
            .I(N__4147));
    Sp12to4 I__823 (
            .O(N__4147),
            .I(N__4144));
    Span12Mux_h I__822 (
            .O(N__4144),
            .I(N__4141));
    Odrv12 I__821 (
            .O(N__4141),
            .I(switch_dn_c));
    InMux I__820 (
            .O(N__4138),
            .I(N__4135));
    LocalMux I__819 (
            .O(N__4135),
            .I(N__4132));
    Odrv12 I__818 (
            .O(N__4132),
            .I(\d2.syncZ0Z_0 ));
    InMux I__817 (
            .O(N__4129),
            .I(N__4125));
    InMux I__816 (
            .O(N__4128),
            .I(N__4122));
    LocalMux I__815 (
            .O(N__4125),
            .I(\d2.syncZ0Z_1 ));
    LocalMux I__814 (
            .O(N__4122),
            .I(\d2.syncZ0Z_1 ));
    InMux I__813 (
            .O(N__4117),
            .I(N__4112));
    CascadeMux I__812 (
            .O(N__4116),
            .I(N__4109));
    CascadeMux I__811 (
            .O(N__4115),
            .I(N__4105));
    LocalMux I__810 (
            .O(N__4112),
            .I(N__4097));
    InMux I__809 (
            .O(N__4109),
            .I(N__4092));
    InMux I__808 (
            .O(N__4108),
            .I(N__4092));
    InMux I__807 (
            .O(N__4105),
            .I(N__4085));
    InMux I__806 (
            .O(N__4104),
            .I(N__4085));
    InMux I__805 (
            .O(N__4103),
            .I(N__4085));
    CascadeMux I__804 (
            .O(N__4102),
            .I(N__4081));
    CascadeMux I__803 (
            .O(N__4101),
            .I(N__4078));
    InMux I__802 (
            .O(N__4100),
            .I(N__4070));
    Span4Mux_h I__801 (
            .O(N__4097),
            .I(N__4063));
    LocalMux I__800 (
            .O(N__4092),
            .I(N__4063));
    LocalMux I__799 (
            .O(N__4085),
            .I(N__4063));
    InMux I__798 (
            .O(N__4084),
            .I(N__4060));
    InMux I__797 (
            .O(N__4081),
            .I(N__4053));
    InMux I__796 (
            .O(N__4078),
            .I(N__4053));
    InMux I__795 (
            .O(N__4077),
            .I(N__4053));
    InMux I__794 (
            .O(N__4076),
            .I(N__4050));
    InMux I__793 (
            .O(N__4075),
            .I(N__4043));
    InMux I__792 (
            .O(N__4074),
            .I(N__4043));
    InMux I__791 (
            .O(N__4073),
            .I(N__4043));
    LocalMux I__790 (
            .O(N__4070),
            .I(d2_state));
    Odrv4 I__789 (
            .O(N__4063),
            .I(d2_state));
    LocalMux I__788 (
            .O(N__4060),
            .I(d2_state));
    LocalMux I__787 (
            .O(N__4053),
            .I(d2_state));
    LocalMux I__786 (
            .O(N__4050),
            .I(d2_state));
    LocalMux I__785 (
            .O(N__4043),
            .I(d2_state));
    IoInMux I__784 (
            .O(N__4030),
            .I(N__4027));
    LocalMux I__783 (
            .O(N__4027),
            .I(N__4024));
    Span4Mux_s1_v I__782 (
            .O(N__4024),
            .I(N__4021));
    Sp12to4 I__781 (
            .O(N__4021),
            .I(N__4018));
    Span12Mux_h I__780 (
            .O(N__4018),
            .I(N__4015));
    Span12Mux_v I__779 (
            .O(N__4015),
            .I(N__4012));
    Odrv12 I__778 (
            .O(N__4012),
            .I(\d2.idle_i ));
    InMux I__777 (
            .O(N__4009),
            .I(N__4005));
    InMux I__776 (
            .O(N__4008),
            .I(N__4001));
    LocalMux I__775 (
            .O(N__4005),
            .I(N__3998));
    InMux I__774 (
            .O(N__4004),
            .I(N__3995));
    LocalMux I__773 (
            .O(N__4001),
            .I(\d1.countZ0Z_1 ));
    Odrv4 I__772 (
            .O(N__3998),
            .I(\d1.countZ0Z_1 ));
    LocalMux I__771 (
            .O(N__3995),
            .I(\d1.countZ0Z_1 ));
    CascadeMux I__770 (
            .O(N__3988),
            .I(N__3985));
    InMux I__769 (
            .O(N__3985),
            .I(N__3980));
    InMux I__768 (
            .O(N__3984),
            .I(N__3973));
    InMux I__767 (
            .O(N__3983),
            .I(N__3973));
    LocalMux I__766 (
            .O(N__3980),
            .I(N__3970));
    InMux I__765 (
            .O(N__3979),
            .I(N__3965));
    InMux I__764 (
            .O(N__3978),
            .I(N__3965));
    LocalMux I__763 (
            .O(N__3973),
            .I(\d1.countZ0Z_0 ));
    Odrv4 I__762 (
            .O(N__3970),
            .I(\d1.countZ0Z_0 ));
    LocalMux I__761 (
            .O(N__3965),
            .I(\d1.countZ0Z_0 ));
    InMux I__760 (
            .O(N__3958),
            .I(N__3954));
    InMux I__759 (
            .O(N__3957),
            .I(N__3951));
    LocalMux I__758 (
            .O(N__3954),
            .I(\d1.countZ0Z_2 ));
    LocalMux I__757 (
            .O(N__3951),
            .I(\d1.countZ0Z_2 ));
    InMux I__756 (
            .O(N__3946),
            .I(\d1.un3_count_cry_1 ));
    InMux I__755 (
            .O(N__3943),
            .I(N__3939));
    InMux I__754 (
            .O(N__3942),
            .I(N__3935));
    LocalMux I__753 (
            .O(N__3939),
            .I(N__3932));
    InMux I__752 (
            .O(N__3938),
            .I(N__3929));
    LocalMux I__751 (
            .O(N__3935),
            .I(\p.countZ0Z_14 ));
    Odrv4 I__750 (
            .O(N__3932),
            .I(\p.countZ0Z_14 ));
    LocalMux I__749 (
            .O(N__3929),
            .I(\p.countZ0Z_14 ));
    InMux I__748 (
            .O(N__3922),
            .I(N__3917));
    InMux I__747 (
            .O(N__3921),
            .I(N__3914));
    InMux I__746 (
            .O(N__3920),
            .I(N__3911));
    LocalMux I__745 (
            .O(N__3917),
            .I(N__3908));
    LocalMux I__744 (
            .O(N__3914),
            .I(\p.countZ0Z_8 ));
    LocalMux I__743 (
            .O(N__3911),
            .I(\p.countZ0Z_8 ));
    Odrv4 I__742 (
            .O(N__3908),
            .I(\p.countZ0Z_8 ));
    InMux I__741 (
            .O(N__3901),
            .I(N__3896));
    CascadeMux I__740 (
            .O(N__3900),
            .I(N__3893));
    InMux I__739 (
            .O(N__3899),
            .I(N__3890));
    LocalMux I__738 (
            .O(N__3896),
            .I(N__3887));
    InMux I__737 (
            .O(N__3893),
            .I(N__3884));
    LocalMux I__736 (
            .O(N__3890),
            .I(\p.countZ0Z_15 ));
    Odrv4 I__735 (
            .O(N__3887),
            .I(\p.countZ0Z_15 ));
    LocalMux I__734 (
            .O(N__3884),
            .I(\p.countZ0Z_15 ));
    InMux I__733 (
            .O(N__3877),
            .I(N__3872));
    InMux I__732 (
            .O(N__3876),
            .I(N__3869));
    InMux I__731 (
            .O(N__3875),
            .I(N__3866));
    LocalMux I__730 (
            .O(N__3872),
            .I(N__3863));
    LocalMux I__729 (
            .O(N__3869),
            .I(\p.countZ0Z_6 ));
    LocalMux I__728 (
            .O(N__3866),
            .I(\p.countZ0Z_6 ));
    Odrv4 I__727 (
            .O(N__3863),
            .I(\p.countZ0Z_6 ));
    InMux I__726 (
            .O(N__3856),
            .I(N__3851));
    InMux I__725 (
            .O(N__3855),
            .I(N__3848));
    InMux I__724 (
            .O(N__3854),
            .I(N__3845));
    LocalMux I__723 (
            .O(N__3851),
            .I(N__3842));
    LocalMux I__722 (
            .O(N__3848),
            .I(\p.countZ0Z_12 ));
    LocalMux I__721 (
            .O(N__3845),
            .I(\p.countZ0Z_12 ));
    Odrv4 I__720 (
            .O(N__3842),
            .I(\p.countZ0Z_12 ));
    InMux I__719 (
            .O(N__3835),
            .I(N__3830));
    InMux I__718 (
            .O(N__3834),
            .I(N__3827));
    InMux I__717 (
            .O(N__3833),
            .I(N__3824));
    LocalMux I__716 (
            .O(N__3830),
            .I(N__3821));
    LocalMux I__715 (
            .O(N__3827),
            .I(\p.countZ0Z_7 ));
    LocalMux I__714 (
            .O(N__3824),
            .I(\p.countZ0Z_7 ));
    Odrv4 I__713 (
            .O(N__3821),
            .I(\p.countZ0Z_7 ));
    CascadeMux I__712 (
            .O(N__3814),
            .I(N__3809));
    InMux I__711 (
            .O(N__3813),
            .I(N__3806));
    InMux I__710 (
            .O(N__3812),
            .I(N__3803));
    InMux I__709 (
            .O(N__3809),
            .I(N__3800));
    LocalMux I__708 (
            .O(N__3806),
            .I(N__3797));
    LocalMux I__707 (
            .O(N__3803),
            .I(\p.countZ0Z_13 ));
    LocalMux I__706 (
            .O(N__3800),
            .I(\p.countZ0Z_13 ));
    Odrv4 I__705 (
            .O(N__3797),
            .I(\p.countZ0Z_13 ));
    InMux I__704 (
            .O(N__3790),
            .I(N__3785));
    InMux I__703 (
            .O(N__3789),
            .I(N__3782));
    InMux I__702 (
            .O(N__3788),
            .I(N__3779));
    LocalMux I__701 (
            .O(N__3785),
            .I(N__3776));
    LocalMux I__700 (
            .O(N__3782),
            .I(\p.countZ0Z_5 ));
    LocalMux I__699 (
            .O(N__3779),
            .I(\p.countZ0Z_5 ));
    Odrv4 I__698 (
            .O(N__3776),
            .I(\p.countZ0Z_5 ));
    InMux I__697 (
            .O(N__3769),
            .I(N__3764));
    InMux I__696 (
            .O(N__3768),
            .I(N__3761));
    InMux I__695 (
            .O(N__3767),
            .I(N__3758));
    LocalMux I__694 (
            .O(N__3764),
            .I(N__3755));
    LocalMux I__693 (
            .O(N__3761),
            .I(\p.countZ0Z_10 ));
    LocalMux I__692 (
            .O(N__3758),
            .I(\p.countZ0Z_10 ));
    Odrv4 I__691 (
            .O(N__3755),
            .I(\p.countZ0Z_10 ));
    InMux I__690 (
            .O(N__3748),
            .I(N__3743));
    InMux I__689 (
            .O(N__3747),
            .I(N__3740));
    InMux I__688 (
            .O(N__3746),
            .I(N__3737));
    LocalMux I__687 (
            .O(N__3743),
            .I(N__3734));
    LocalMux I__686 (
            .O(N__3740),
            .I(\p.countZ0Z_9 ));
    LocalMux I__685 (
            .O(N__3737),
            .I(\p.countZ0Z_9 ));
    Odrv4 I__684 (
            .O(N__3734),
            .I(\p.countZ0Z_9 ));
    CascadeMux I__683 (
            .O(N__3727),
            .I(N__3722));
    InMux I__682 (
            .O(N__3726),
            .I(N__3719));
    InMux I__681 (
            .O(N__3725),
            .I(N__3716));
    InMux I__680 (
            .O(N__3722),
            .I(N__3713));
    LocalMux I__679 (
            .O(N__3719),
            .I(N__3710));
    LocalMux I__678 (
            .O(N__3716),
            .I(\p.countZ0Z_11 ));
    LocalMux I__677 (
            .O(N__3713),
            .I(\p.countZ0Z_11 ));
    Odrv4 I__676 (
            .O(N__3710),
            .I(\p.countZ0Z_11 ));
    InMux I__675 (
            .O(N__3703),
            .I(N__3698));
    InMux I__674 (
            .O(N__3702),
            .I(N__3695));
    InMux I__673 (
            .O(N__3701),
            .I(N__3692));
    LocalMux I__672 (
            .O(N__3698),
            .I(N__3689));
    LocalMux I__671 (
            .O(N__3695),
            .I(\p.countZ0Z_4 ));
    LocalMux I__670 (
            .O(N__3692),
            .I(\p.countZ0Z_4 ));
    Odrv4 I__669 (
            .O(N__3689),
            .I(\p.countZ0Z_4 ));
    InMux I__668 (
            .O(N__3682),
            .I(N__3679));
    LocalMux I__667 (
            .O(N__3679),
            .I(\p.count10_11 ));
    InMux I__666 (
            .O(N__3676),
            .I(N__3673));
    LocalMux I__665 (
            .O(N__3673),
            .I(\p.count10_10 ));
    CascadeMux I__664 (
            .O(N__3670),
            .I(\p.count10_8_cascade_ ));
    InMux I__663 (
            .O(N__3667),
            .I(N__3658));
    InMux I__662 (
            .O(N__3666),
            .I(N__3658));
    InMux I__661 (
            .O(N__3665),
            .I(N__3655));
    InMux I__660 (
            .O(N__3664),
            .I(N__3650));
    InMux I__659 (
            .O(N__3663),
            .I(N__3650));
    LocalMux I__658 (
            .O(N__3658),
            .I(\p.count10 ));
    LocalMux I__657 (
            .O(N__3655),
            .I(\p.count10 ));
    LocalMux I__656 (
            .O(N__3650),
            .I(\p.count10 ));
    InMux I__655 (
            .O(N__3643),
            .I(N__3638));
    InMux I__654 (
            .O(N__3642),
            .I(N__3635));
    InMux I__653 (
            .O(N__3641),
            .I(N__3632));
    LocalMux I__652 (
            .O(N__3638),
            .I(N__3629));
    LocalMux I__651 (
            .O(N__3635),
            .I(\p.countZ0Z_3 ));
    LocalMux I__650 (
            .O(N__3632),
            .I(\p.countZ0Z_3 ));
    Odrv4 I__649 (
            .O(N__3629),
            .I(\p.countZ0Z_3 ));
    InMux I__648 (
            .O(N__3622),
            .I(N__3617));
    InMux I__647 (
            .O(N__3621),
            .I(N__3614));
    InMux I__646 (
            .O(N__3620),
            .I(N__3611));
    LocalMux I__645 (
            .O(N__3617),
            .I(N__3608));
    LocalMux I__644 (
            .O(N__3614),
            .I(\p.countZ0Z_2 ));
    LocalMux I__643 (
            .O(N__3611),
            .I(\p.countZ0Z_2 ));
    Odrv4 I__642 (
            .O(N__3608),
            .I(\p.countZ0Z_2 ));
    InMux I__641 (
            .O(N__3601),
            .I(N__3598));
    LocalMux I__640 (
            .O(N__3598),
            .I(\p.count10_9 ));
    InMux I__639 (
            .O(N__3595),
            .I(N__3592));
    LocalMux I__638 (
            .O(N__3592),
            .I(N__3589));
    Span4Mux_v I__637 (
            .O(N__3589),
            .I(N__3586));
    Odrv4 I__636 (
            .O(N__3586),
            .I(\d2.trans_up_1_11 ));
    InMux I__635 (
            .O(N__3583),
            .I(N__3580));
    LocalMux I__634 (
            .O(N__3580),
            .I(N__3577));
    Span4Mux_v I__633 (
            .O(N__3577),
            .I(N__3574));
    Odrv4 I__632 (
            .O(N__3574),
            .I(\d2.trans_up_1_10 ));
    InMux I__631 (
            .O(N__3571),
            .I(N__3568));
    LocalMux I__630 (
            .O(N__3568),
            .I(\d1.trans_up_1_11 ));
    CascadeMux I__629 (
            .O(N__3565),
            .I(\d1.trans_up_1_13_sx_cascade_ ));
    InMux I__628 (
            .O(N__3562),
            .I(N__3559));
    LocalMux I__627 (
            .O(N__3559),
            .I(\d1.trans_up_1_14 ));
    CascadeMux I__626 (
            .O(N__3556),
            .I(\d1.trans_up_1_13_cascade_ ));
    InMux I__625 (
            .O(N__3553),
            .I(N__3549));
    InMux I__624 (
            .O(N__3552),
            .I(N__3546));
    LocalMux I__623 (
            .O(N__3549),
            .I(\d1.trans_up_1_12 ));
    LocalMux I__622 (
            .O(N__3546),
            .I(\d1.trans_up_1_12 ));
    InMux I__621 (
            .O(N__3541),
            .I(N__3538));
    LocalMux I__620 (
            .O(N__3538),
            .I(\d1.trans_up_1_9 ));
    InMux I__619 (
            .O(N__3535),
            .I(N__3532));
    LocalMux I__618 (
            .O(N__3532),
            .I(\d1.trans_up_sx ));
    InMux I__617 (
            .O(N__3529),
            .I(N__3517));
    InMux I__616 (
            .O(N__3528),
            .I(N__3517));
    InMux I__615 (
            .O(N__3527),
            .I(N__3517));
    InMux I__614 (
            .O(N__3526),
            .I(N__3517));
    LocalMux I__613 (
            .O(N__3517),
            .I(\d1.stateZ0 ));
    CascadeMux I__612 (
            .O(N__3514),
            .I(N__3510));
    InMux I__611 (
            .O(N__3513),
            .I(N__3507));
    InMux I__610 (
            .O(N__3510),
            .I(N__3504));
    LocalMux I__609 (
            .O(N__3507),
            .I(\d1.syncZ0Z_1 ));
    LocalMux I__608 (
            .O(N__3504),
            .I(\d1.syncZ0Z_1 ));
    IoInMux I__607 (
            .O(N__3499),
            .I(N__3496));
    LocalMux I__606 (
            .O(N__3496),
            .I(N__3493));
    Span12Mux_s8_h I__605 (
            .O(N__3493),
            .I(N__3490));
    Odrv12 I__604 (
            .O(N__3490),
            .I(\d1.idle_i ));
    CascadeMux I__603 (
            .O(N__3487),
            .I(N__3484));
    InMux I__602 (
            .O(N__3484),
            .I(N__3481));
    LocalMux I__601 (
            .O(N__3481),
            .I(state_RNIU5D07));
    InMux I__600 (
            .O(N__3478),
            .I(N__3475));
    LocalMux I__599 (
            .O(N__3475),
            .I(state_RNIPC4P3_1));
    InMux I__598 (
            .O(N__3472),
            .I(N__3469));
    LocalMux I__597 (
            .O(N__3469),
            .I(state_RNIPC4P3_8));
    InMux I__596 (
            .O(N__3466),
            .I(N__3448));
    InMux I__595 (
            .O(N__3465),
            .I(N__3448));
    InMux I__594 (
            .O(N__3464),
            .I(N__3448));
    InMux I__593 (
            .O(N__3463),
            .I(N__3441));
    InMux I__592 (
            .O(N__3462),
            .I(N__3441));
    InMux I__591 (
            .O(N__3461),
            .I(N__3441));
    InMux I__590 (
            .O(N__3460),
            .I(N__3438));
    InMux I__589 (
            .O(N__3459),
            .I(N__3431));
    InMux I__588 (
            .O(N__3458),
            .I(N__3431));
    InMux I__587 (
            .O(N__3457),
            .I(N__3431));
    InMux I__586 (
            .O(N__3456),
            .I(N__3426));
    InMux I__585 (
            .O(N__3455),
            .I(N__3426));
    LocalMux I__584 (
            .O(N__3448),
            .I(d2_trans_up_1));
    LocalMux I__583 (
            .O(N__3441),
            .I(d2_trans_up_1));
    LocalMux I__582 (
            .O(N__3438),
            .I(d2_trans_up_1));
    LocalMux I__581 (
            .O(N__3431),
            .I(d2_trans_up_1));
    LocalMux I__580 (
            .O(N__3426),
            .I(d2_trans_up_1));
    InMux I__579 (
            .O(N__3415),
            .I(N__3412));
    LocalMux I__578 (
            .O(N__3412),
            .I(state_RNIPC4P3_5));
    CascadeMux I__577 (
            .O(N__3409),
            .I(\d1.count_RNI2PCEZ0Z_3_cascade_ ));
    CascadeMux I__576 (
            .O(N__3406),
            .I(\d1.trans_up_1_14_cascade_ ));
    CascadeMux I__575 (
            .O(N__3403),
            .I(N__3400));
    InMux I__574 (
            .O(N__3400),
            .I(N__3391));
    InMux I__573 (
            .O(N__3399),
            .I(N__3391));
    InMux I__572 (
            .O(N__3398),
            .I(N__3391));
    LocalMux I__571 (
            .O(N__3391),
            .I(s_up));
    CascadeMux I__570 (
            .O(N__3388),
            .I(s_up_cascade_));
    InMux I__569 (
            .O(N__3385),
            .I(N__3378));
    InMux I__568 (
            .O(N__3384),
            .I(N__3378));
    InMux I__567 (
            .O(N__3383),
            .I(N__3375));
    LocalMux I__566 (
            .O(N__3378),
            .I(s_dn_i));
    LocalMux I__565 (
            .O(N__3375),
            .I(s_dn_i));
    CascadeMux I__564 (
            .O(N__3370),
            .I(N__3367));
    InMux I__563 (
            .O(N__3367),
            .I(N__3364));
    LocalMux I__562 (
            .O(N__3364),
            .I(state_RNIU5D07_0));
    InMux I__561 (
            .O(N__3361),
            .I(N__3358));
    LocalMux I__560 (
            .O(N__3358),
            .I(state_RNIPC4P3_0));
    InMux I__559 (
            .O(N__3355),
            .I(N__3352));
    LocalMux I__558 (
            .O(N__3352),
            .I(state_RNIPC4P3_2));
    CascadeMux I__557 (
            .O(N__3349),
            .I(\d2.trans_up_1_12_cascade_ ));
    CascadeMux I__556 (
            .O(N__3346),
            .I(\d2.trans_up_1_sx_cascade_ ));
    CascadeMux I__555 (
            .O(N__3343),
            .I(d2_trans_up_1_cascade_));
    CascadeMux I__554 (
            .O(N__3340),
            .I(N__3337));
    InMux I__553 (
            .O(N__3337),
            .I(N__3332));
    InMux I__552 (
            .O(N__3336),
            .I(N__3326));
    InMux I__551 (
            .O(N__3335),
            .I(N__3326));
    LocalMux I__550 (
            .O(N__3332),
            .I(N__3323));
    InMux I__549 (
            .O(N__3331),
            .I(N__3320));
    LocalMux I__548 (
            .O(N__3326),
            .I(N__3315));
    Span4Mux_h I__547 (
            .O(N__3323),
            .I(N__3315));
    LocalMux I__546 (
            .O(N__3320),
            .I(pulse_lenZ0Z_2));
    Odrv4 I__545 (
            .O(N__3315),
            .I(pulse_lenZ0Z_2));
    CascadeMux I__544 (
            .O(N__3310),
            .I(s_dn_i_cascade_));
    CascadeMux I__543 (
            .O(N__3307),
            .I(N__3304));
    InMux I__542 (
            .O(N__3304),
            .I(N__3301));
    LocalMux I__541 (
            .O(N__3301),
            .I(un1_pulse_len_cry_2_c_RNOZ0));
    InMux I__540 (
            .O(N__3298),
            .I(N__3295));
    LocalMux I__539 (
            .O(N__3295),
            .I(state_RNIPC4P3_3));
    InMux I__538 (
            .O(N__3292),
            .I(\p.count_1_cry_7 ));
    InMux I__537 (
            .O(N__3289),
            .I(bfn_7_13_0_));
    InMux I__536 (
            .O(N__3286),
            .I(\p.count_1_cry_9 ));
    InMux I__535 (
            .O(N__3283),
            .I(\p.count_1_cry_10 ));
    InMux I__534 (
            .O(N__3280),
            .I(\p.count_1_cry_11 ));
    InMux I__533 (
            .O(N__3277),
            .I(\p.count_1_cry_12 ));
    InMux I__532 (
            .O(N__3274),
            .I(\p.count_1_cry_13 ));
    InMux I__531 (
            .O(N__3271),
            .I(\p.count_1_cry_14 ));
    CascadeMux I__530 (
            .O(N__3268),
            .I(N__3265));
    InMux I__529 (
            .O(N__3265),
            .I(N__3261));
    CascadeMux I__528 (
            .O(N__3264),
            .I(N__3258));
    LocalMux I__527 (
            .O(N__3261),
            .I(N__3255));
    InMux I__526 (
            .O(N__3258),
            .I(N__3252));
    Span4Mux_h I__525 (
            .O(N__3255),
            .I(N__3249));
    LocalMux I__524 (
            .O(N__3252),
            .I(pulse_lenZ0Z_15));
    Odrv4 I__523 (
            .O(N__3249),
            .I(pulse_lenZ0Z_15));
    InMux I__522 (
            .O(N__3244),
            .I(N__3241));
    LocalMux I__521 (
            .O(N__3241),
            .I(\p.count_i_15 ));
    InMux I__520 (
            .O(N__3238),
            .I(\p.CONTROL_PIN_2 ));
    IoInMux I__519 (
            .O(N__3235),
            .I(N__3232));
    LocalMux I__518 (
            .O(N__3232),
            .I(N__3229));
    IoSpan4Mux I__517 (
            .O(N__3229),
            .I(N__3226));
    Sp12to4 I__516 (
            .O(N__3226),
            .I(N__3223));
    Span12Mux_h I__515 (
            .O(N__3223),
            .I(N__3220));
    Span12Mux_v I__514 (
            .O(N__3220),
            .I(N__3217));
    Odrv12 I__513 (
            .O(N__3217),
            .I(CONTROL_PIN_c));
    InMux I__512 (
            .O(N__3214),
            .I(\p.count_1_cry_1 ));
    InMux I__511 (
            .O(N__3211),
            .I(\p.count_1_cry_2 ));
    InMux I__510 (
            .O(N__3208),
            .I(\p.count_1_cry_3 ));
    InMux I__509 (
            .O(N__3205),
            .I(\p.count_1_cry_4 ));
    InMux I__508 (
            .O(N__3202),
            .I(\p.count_1_cry_5 ));
    InMux I__507 (
            .O(N__3199),
            .I(\p.count_1_cry_6 ));
    CascadeMux I__506 (
            .O(N__3196),
            .I(N__3193));
    InMux I__505 (
            .O(N__3193),
            .I(N__3189));
    CascadeMux I__504 (
            .O(N__3192),
            .I(N__3186));
    LocalMux I__503 (
            .O(N__3189),
            .I(N__3183));
    InMux I__502 (
            .O(N__3186),
            .I(N__3180));
    Span4Mux_h I__501 (
            .O(N__3183),
            .I(N__3177));
    LocalMux I__500 (
            .O(N__3180),
            .I(pulse_lenZ0Z_7));
    Odrv4 I__499 (
            .O(N__3177),
            .I(pulse_lenZ0Z_7));
    InMux I__498 (
            .O(N__3172),
            .I(N__3169));
    LocalMux I__497 (
            .O(N__3169),
            .I(\p.count_i_7 ));
    CascadeMux I__496 (
            .O(N__3166),
            .I(N__3162));
    CascadeMux I__495 (
            .O(N__3165),
            .I(N__3159));
    InMux I__494 (
            .O(N__3162),
            .I(N__3156));
    InMux I__493 (
            .O(N__3159),
            .I(N__3153));
    LocalMux I__492 (
            .O(N__3156),
            .I(N__3150));
    LocalMux I__491 (
            .O(N__3153),
            .I(N__3145));
    Span4Mux_h I__490 (
            .O(N__3150),
            .I(N__3145));
    Odrv4 I__489 (
            .O(N__3145),
            .I(pulse_lenZ0Z_8));
    InMux I__488 (
            .O(N__3142),
            .I(N__3139));
    LocalMux I__487 (
            .O(N__3139),
            .I(\p.count_i_8 ));
    CascadeMux I__486 (
            .O(N__3136),
            .I(N__3132));
    InMux I__485 (
            .O(N__3135),
            .I(N__3129));
    InMux I__484 (
            .O(N__3132),
            .I(N__3126));
    LocalMux I__483 (
            .O(N__3129),
            .I(N__3123));
    LocalMux I__482 (
            .O(N__3126),
            .I(pulse_lenZ0Z_9));
    Odrv4 I__481 (
            .O(N__3123),
            .I(pulse_lenZ0Z_9));
    CascadeMux I__480 (
            .O(N__3118),
            .I(N__3115));
    InMux I__479 (
            .O(N__3115),
            .I(N__3112));
    LocalMux I__478 (
            .O(N__3112),
            .I(\p.count_i_9 ));
    CascadeMux I__477 (
            .O(N__3109),
            .I(N__3105));
    CascadeMux I__476 (
            .O(N__3108),
            .I(N__3102));
    InMux I__475 (
            .O(N__3105),
            .I(N__3099));
    InMux I__474 (
            .O(N__3102),
            .I(N__3096));
    LocalMux I__473 (
            .O(N__3099),
            .I(N__3093));
    LocalMux I__472 (
            .O(N__3096),
            .I(pulse_lenZ0Z_10));
    Odrv4 I__471 (
            .O(N__3093),
            .I(pulse_lenZ0Z_10));
    InMux I__470 (
            .O(N__3088),
            .I(N__3085));
    LocalMux I__469 (
            .O(N__3085),
            .I(\p.count_i_10 ));
    CascadeMux I__468 (
            .O(N__3082),
            .I(N__3079));
    InMux I__467 (
            .O(N__3079),
            .I(N__3075));
    CascadeMux I__466 (
            .O(N__3078),
            .I(N__3072));
    LocalMux I__465 (
            .O(N__3075),
            .I(N__3069));
    InMux I__464 (
            .O(N__3072),
            .I(N__3066));
    Span4Mux_h I__463 (
            .O(N__3069),
            .I(N__3063));
    LocalMux I__462 (
            .O(N__3066),
            .I(pulse_lenZ0Z_11));
    Odrv4 I__461 (
            .O(N__3063),
            .I(pulse_lenZ0Z_11));
    InMux I__460 (
            .O(N__3058),
            .I(N__3055));
    LocalMux I__459 (
            .O(N__3055),
            .I(\p.count_i_11 ));
    CascadeMux I__458 (
            .O(N__3052),
            .I(N__3048));
    CascadeMux I__457 (
            .O(N__3051),
            .I(N__3045));
    InMux I__456 (
            .O(N__3048),
            .I(N__3042));
    InMux I__455 (
            .O(N__3045),
            .I(N__3039));
    LocalMux I__454 (
            .O(N__3042),
            .I(N__3036));
    LocalMux I__453 (
            .O(N__3039),
            .I(pulse_lenZ0Z_12));
    Odrv4 I__452 (
            .O(N__3036),
            .I(pulse_lenZ0Z_12));
    InMux I__451 (
            .O(N__3031),
            .I(N__3028));
    LocalMux I__450 (
            .O(N__3028),
            .I(\p.count_i_12 ));
    CascadeMux I__449 (
            .O(N__3025),
            .I(N__3021));
    CascadeMux I__448 (
            .O(N__3024),
            .I(N__3018));
    InMux I__447 (
            .O(N__3021),
            .I(N__3015));
    InMux I__446 (
            .O(N__3018),
            .I(N__3012));
    LocalMux I__445 (
            .O(N__3015),
            .I(N__3009));
    LocalMux I__444 (
            .O(N__3012),
            .I(pulse_lenZ0Z_13));
    Odrv4 I__443 (
            .O(N__3009),
            .I(pulse_lenZ0Z_13));
    InMux I__442 (
            .O(N__3004),
            .I(N__3001));
    LocalMux I__441 (
            .O(N__3001),
            .I(\p.count_i_13 ));
    CascadeMux I__440 (
            .O(N__2998),
            .I(N__2994));
    CascadeMux I__439 (
            .O(N__2997),
            .I(N__2991));
    InMux I__438 (
            .O(N__2994),
            .I(N__2988));
    InMux I__437 (
            .O(N__2991),
            .I(N__2985));
    LocalMux I__436 (
            .O(N__2988),
            .I(N__2982));
    LocalMux I__435 (
            .O(N__2985),
            .I(pulse_lenZ0Z_14));
    Odrv4 I__434 (
            .O(N__2982),
            .I(pulse_lenZ0Z_14));
    InMux I__433 (
            .O(N__2977),
            .I(N__2974));
    LocalMux I__432 (
            .O(N__2974),
            .I(\p.count_i_14 ));
    InMux I__431 (
            .O(N__2971),
            .I(un1_pulse_len_cry_14));
    InMux I__430 (
            .O(N__2968),
            .I(N__2965));
    LocalMux I__429 (
            .O(N__2965),
            .I(state_RNIPC4P3_4));
    InMux I__428 (
            .O(N__2962),
            .I(N__2959));
    LocalMux I__427 (
            .O(N__2959),
            .I(state_RNIPC4P3_7));
    InMux I__426 (
            .O(N__2956),
            .I(N__2953));
    LocalMux I__425 (
            .O(N__2953),
            .I(\p.count_i_2 ));
    CascadeMux I__424 (
            .O(N__2950),
            .I(N__2947));
    InMux I__423 (
            .O(N__2947),
            .I(N__2943));
    CascadeMux I__422 (
            .O(N__2946),
            .I(N__2940));
    LocalMux I__421 (
            .O(N__2943),
            .I(N__2937));
    InMux I__420 (
            .O(N__2940),
            .I(N__2934));
    Span4Mux_h I__419 (
            .O(N__2937),
            .I(N__2931));
    LocalMux I__418 (
            .O(N__2934),
            .I(pulse_lenZ0Z_3));
    Odrv4 I__417 (
            .O(N__2931),
            .I(pulse_lenZ0Z_3));
    InMux I__416 (
            .O(N__2926),
            .I(N__2923));
    LocalMux I__415 (
            .O(N__2923),
            .I(\p.count_i_3 ));
    CascadeMux I__414 (
            .O(N__2920),
            .I(N__2916));
    CascadeMux I__413 (
            .O(N__2919),
            .I(N__2913));
    InMux I__412 (
            .O(N__2916),
            .I(N__2910));
    InMux I__411 (
            .O(N__2913),
            .I(N__2907));
    LocalMux I__410 (
            .O(N__2910),
            .I(N__2904));
    LocalMux I__409 (
            .O(N__2907),
            .I(pulse_lenZ0Z_4));
    Odrv4 I__408 (
            .O(N__2904),
            .I(pulse_lenZ0Z_4));
    InMux I__407 (
            .O(N__2899),
            .I(N__2896));
    LocalMux I__406 (
            .O(N__2896),
            .I(\p.count_i_4 ));
    CascadeMux I__405 (
            .O(N__2893),
            .I(N__2890));
    InMux I__404 (
            .O(N__2890),
            .I(N__2887));
    LocalMux I__403 (
            .O(N__2887),
            .I(N__2883));
    InMux I__402 (
            .O(N__2886),
            .I(N__2880));
    Span4Mux_v I__401 (
            .O(N__2883),
            .I(N__2877));
    LocalMux I__400 (
            .O(N__2880),
            .I(pulse_lenZ0Z_5));
    Odrv4 I__399 (
            .O(N__2877),
            .I(pulse_lenZ0Z_5));
    InMux I__398 (
            .O(N__2872),
            .I(N__2869));
    LocalMux I__397 (
            .O(N__2869),
            .I(\p.count_i_5 ));
    CascadeMux I__396 (
            .O(N__2866),
            .I(N__2863));
    InMux I__395 (
            .O(N__2863),
            .I(N__2859));
    InMux I__394 (
            .O(N__2862),
            .I(N__2856));
    LocalMux I__393 (
            .O(N__2859),
            .I(N__2853));
    LocalMux I__392 (
            .O(N__2856),
            .I(pulse_lenZ0Z_6));
    Odrv4 I__391 (
            .O(N__2853),
            .I(pulse_lenZ0Z_6));
    InMux I__390 (
            .O(N__2848),
            .I(N__2845));
    LocalMux I__389 (
            .O(N__2845),
            .I(\p.count_i_6 ));
    InMux I__388 (
            .O(N__2842),
            .I(un1_pulse_len_cry_5));
    InMux I__387 (
            .O(N__2839),
            .I(un1_pulse_len_cry_6));
    InMux I__386 (
            .O(N__2836),
            .I(N__2833));
    LocalMux I__385 (
            .O(N__2833),
            .I(state_RNIPC4P3_6));
    InMux I__384 (
            .O(N__2830),
            .I(un1_pulse_len_cry_7));
    InMux I__383 (
            .O(N__2827),
            .I(un1_pulse_len_cry_8));
    InMux I__382 (
            .O(N__2824),
            .I(bfn_7_9_0_));
    InMux I__381 (
            .O(N__2821),
            .I(un1_pulse_len_cry_10));
    InMux I__380 (
            .O(N__2818),
            .I(un1_pulse_len_cry_11));
    InMux I__379 (
            .O(N__2815),
            .I(un1_pulse_len_cry_12));
    InMux I__378 (
            .O(N__2812),
            .I(un1_pulse_len_cry_13));
    InMux I__377 (
            .O(N__2809),
            .I(N__2806));
    LocalMux I__376 (
            .O(N__2806),
            .I(\p.prescaler_1_cry_5_THRU_CO ));
    CascadeMux I__375 (
            .O(N__2803),
            .I(N__2798));
    CascadeMux I__374 (
            .O(N__2802),
            .I(N__2795));
    InMux I__373 (
            .O(N__2801),
            .I(N__2792));
    InMux I__372 (
            .O(N__2798),
            .I(N__2787));
    InMux I__371 (
            .O(N__2795),
            .I(N__2787));
    LocalMux I__370 (
            .O(N__2792),
            .I(\p.prescalerZ0Z_6 ));
    LocalMux I__369 (
            .O(N__2787),
            .I(\p.prescalerZ0Z_6 ));
    InMux I__368 (
            .O(N__2782),
            .I(N__2779));
    LocalMux I__367 (
            .O(N__2779),
            .I(\p.prescaler_1_cry_4_THRU_CO ));
    InMux I__366 (
            .O(N__2776),
            .I(N__2771));
    InMux I__365 (
            .O(N__2775),
            .I(N__2766));
    InMux I__364 (
            .O(N__2774),
            .I(N__2766));
    LocalMux I__363 (
            .O(N__2771),
            .I(\p.prescalerZ0Z_5 ));
    LocalMux I__362 (
            .O(N__2766),
            .I(\p.prescalerZ0Z_5 ));
    InMux I__361 (
            .O(N__2761),
            .I(N__2755));
    InMux I__360 (
            .O(N__2760),
            .I(N__2748));
    InMux I__359 (
            .O(N__2759),
            .I(N__2748));
    InMux I__358 (
            .O(N__2758),
            .I(N__2748));
    LocalMux I__357 (
            .O(N__2755),
            .I(\p.prescalerZ0Z_0 ));
    LocalMux I__356 (
            .O(N__2748),
            .I(\p.prescalerZ0Z_0 ));
    CascadeMux I__355 (
            .O(N__2743),
            .I(N__2740));
    InMux I__354 (
            .O(N__2740),
            .I(N__2735));
    InMux I__353 (
            .O(N__2739),
            .I(N__2730));
    InMux I__352 (
            .O(N__2738),
            .I(N__2730));
    LocalMux I__351 (
            .O(N__2735),
            .I(\p.prescalerZ0Z_1 ));
    LocalMux I__350 (
            .O(N__2730),
            .I(\p.prescalerZ0Z_1 ));
    InMux I__349 (
            .O(N__2725),
            .I(N__2722));
    LocalMux I__348 (
            .O(N__2722),
            .I(state_RNIPC4P3));
    InMux I__347 (
            .O(N__2719),
            .I(un1_pulse_len_cry_2));
    InMux I__346 (
            .O(N__2716),
            .I(un1_pulse_len_cry_3));
    InMux I__345 (
            .O(N__2713),
            .I(un1_pulse_len_cry_4));
    InMux I__344 (
            .O(N__2710),
            .I(N__2706));
    InMux I__343 (
            .O(N__2709),
            .I(N__2703));
    LocalMux I__342 (
            .O(N__2706),
            .I(\p.prescalerZ0Z_20 ));
    LocalMux I__341 (
            .O(N__2703),
            .I(\p.prescalerZ0Z_20 ));
    InMux I__340 (
            .O(N__2698),
            .I(\p.prescaler_1_cry_19 ));
    InMux I__339 (
            .O(N__2695),
            .I(N__2691));
    InMux I__338 (
            .O(N__2694),
            .I(N__2688));
    LocalMux I__337 (
            .O(N__2691),
            .I(\p.prescalerZ0Z_21 ));
    LocalMux I__336 (
            .O(N__2688),
            .I(\p.prescalerZ0Z_21 ));
    InMux I__335 (
            .O(N__2683),
            .I(\p.prescaler_1_cry_20 ));
    CascadeMux I__334 (
            .O(N__2680),
            .I(N__2676));
    InMux I__333 (
            .O(N__2679),
            .I(N__2673));
    InMux I__332 (
            .O(N__2676),
            .I(N__2670));
    LocalMux I__331 (
            .O(N__2673),
            .I(\p.prescalerZ0Z_22 ));
    LocalMux I__330 (
            .O(N__2670),
            .I(\p.prescalerZ0Z_22 ));
    InMux I__329 (
            .O(N__2665),
            .I(\p.prescaler_1_cry_21 ));
    CascadeMux I__328 (
            .O(N__2662),
            .I(N__2658));
    InMux I__327 (
            .O(N__2661),
            .I(N__2655));
    InMux I__326 (
            .O(N__2658),
            .I(N__2652));
    LocalMux I__325 (
            .O(N__2655),
            .I(\p.prescalerZ0Z_23 ));
    LocalMux I__324 (
            .O(N__2652),
            .I(\p.prescalerZ0Z_23 ));
    InMux I__323 (
            .O(N__2647),
            .I(\p.prescaler_1_cry_22 ));
    CascadeMux I__322 (
            .O(N__2644),
            .I(N__2641));
    InMux I__321 (
            .O(N__2641),
            .I(N__2637));
    InMux I__320 (
            .O(N__2640),
            .I(N__2634));
    LocalMux I__319 (
            .O(N__2637),
            .I(N__2631));
    LocalMux I__318 (
            .O(N__2634),
            .I(\p.prescalerZ0Z_24 ));
    Odrv4 I__317 (
            .O(N__2631),
            .I(\p.prescalerZ0Z_24 ));
    InMux I__316 (
            .O(N__2626),
            .I(\p.prescaler_1_cry_23 ));
    CascadeMux I__315 (
            .O(N__2623),
            .I(N__2620));
    InMux I__314 (
            .O(N__2620),
            .I(N__2616));
    InMux I__313 (
            .O(N__2619),
            .I(N__2613));
    LocalMux I__312 (
            .O(N__2616),
            .I(N__2610));
    LocalMux I__311 (
            .O(N__2613),
            .I(\p.prescalerZ0Z_25 ));
    Odrv4 I__310 (
            .O(N__2610),
            .I(\p.prescalerZ0Z_25 ));
    InMux I__309 (
            .O(N__2605),
            .I(bfn_2_14_0_));
    InMux I__308 (
            .O(N__2602),
            .I(\p.prescaler_1_cry_25 ));
    CascadeMux I__307 (
            .O(N__2599),
            .I(N__2595));
    InMux I__306 (
            .O(N__2598),
            .I(N__2592));
    InMux I__305 (
            .O(N__2595),
            .I(N__2589));
    LocalMux I__304 (
            .O(N__2592),
            .I(\p.prescalerZ0Z_26 ));
    LocalMux I__303 (
            .O(N__2589),
            .I(\p.prescalerZ0Z_26 ));
    InMux I__302 (
            .O(N__2584),
            .I(N__2581));
    LocalMux I__301 (
            .O(N__2581),
            .I(N__2578));
    Odrv4 I__300 (
            .O(N__2578),
            .I(\p.prescaler12_0_and ));
    InMux I__299 (
            .O(N__2575),
            .I(N__2571));
    InMux I__298 (
            .O(N__2574),
            .I(N__2568));
    LocalMux I__297 (
            .O(N__2571),
            .I(\p.prescalerZ0Z_12 ));
    LocalMux I__296 (
            .O(N__2568),
            .I(\p.prescalerZ0Z_12 ));
    InMux I__295 (
            .O(N__2563),
            .I(\p.prescaler_1_cry_11 ));
    InMux I__294 (
            .O(N__2560),
            .I(N__2556));
    InMux I__293 (
            .O(N__2559),
            .I(N__2553));
    LocalMux I__292 (
            .O(N__2556),
            .I(\p.prescalerZ0Z_13 ));
    LocalMux I__291 (
            .O(N__2553),
            .I(\p.prescalerZ0Z_13 ));
    InMux I__290 (
            .O(N__2548),
            .I(\p.prescaler_1_cry_12 ));
    InMux I__289 (
            .O(N__2545),
            .I(N__2541));
    InMux I__288 (
            .O(N__2544),
            .I(N__2538));
    LocalMux I__287 (
            .O(N__2541),
            .I(\p.prescalerZ0Z_14 ));
    LocalMux I__286 (
            .O(N__2538),
            .I(\p.prescalerZ0Z_14 ));
    InMux I__285 (
            .O(N__2533),
            .I(\p.prescaler_1_cry_13 ));
    InMux I__284 (
            .O(N__2530),
            .I(N__2526));
    InMux I__283 (
            .O(N__2529),
            .I(N__2523));
    LocalMux I__282 (
            .O(N__2526),
            .I(\p.prescalerZ0Z_15 ));
    LocalMux I__281 (
            .O(N__2523),
            .I(\p.prescalerZ0Z_15 ));
    InMux I__280 (
            .O(N__2518),
            .I(\p.prescaler_1_cry_14 ));
    InMux I__279 (
            .O(N__2515),
            .I(N__2511));
    InMux I__278 (
            .O(N__2514),
            .I(N__2508));
    LocalMux I__277 (
            .O(N__2511),
            .I(\p.prescalerZ0Z_16 ));
    LocalMux I__276 (
            .O(N__2508),
            .I(\p.prescalerZ0Z_16 ));
    InMux I__275 (
            .O(N__2503),
            .I(\p.prescaler_1_cry_15 ));
    InMux I__274 (
            .O(N__2500),
            .I(N__2496));
    InMux I__273 (
            .O(N__2499),
            .I(N__2493));
    LocalMux I__272 (
            .O(N__2496),
            .I(\p.prescalerZ0Z_17 ));
    LocalMux I__271 (
            .O(N__2493),
            .I(\p.prescalerZ0Z_17 ));
    InMux I__270 (
            .O(N__2488),
            .I(bfn_2_13_0_));
    InMux I__269 (
            .O(N__2485),
            .I(N__2481));
    InMux I__268 (
            .O(N__2484),
            .I(N__2478));
    LocalMux I__267 (
            .O(N__2481),
            .I(N__2475));
    LocalMux I__266 (
            .O(N__2478),
            .I(\p.prescalerZ0Z_18 ));
    Odrv4 I__265 (
            .O(N__2475),
            .I(\p.prescalerZ0Z_18 ));
    InMux I__264 (
            .O(N__2470),
            .I(\p.prescaler_1_cry_17 ));
    InMux I__263 (
            .O(N__2467),
            .I(N__2463));
    InMux I__262 (
            .O(N__2466),
            .I(N__2460));
    LocalMux I__261 (
            .O(N__2463),
            .I(\p.prescalerZ0Z_19 ));
    LocalMux I__260 (
            .O(N__2460),
            .I(\p.prescalerZ0Z_19 ));
    InMux I__259 (
            .O(N__2455),
            .I(\p.prescaler_1_cry_18 ));
    InMux I__258 (
            .O(N__2452),
            .I(N__2448));
    InMux I__257 (
            .O(N__2451),
            .I(N__2445));
    LocalMux I__256 (
            .O(N__2448),
            .I(\p.prescalerZ0Z_3 ));
    LocalMux I__255 (
            .O(N__2445),
            .I(\p.prescalerZ0Z_3 ));
    InMux I__254 (
            .O(N__2440),
            .I(\p.prescaler_1_cry_2 ));
    InMux I__253 (
            .O(N__2437),
            .I(N__2433));
    InMux I__252 (
            .O(N__2436),
            .I(N__2430));
    LocalMux I__251 (
            .O(N__2433),
            .I(\p.prescalerZ0Z_4 ));
    LocalMux I__250 (
            .O(N__2430),
            .I(\p.prescalerZ0Z_4 ));
    InMux I__249 (
            .O(N__2425),
            .I(\p.prescaler_1_cry_3 ));
    InMux I__248 (
            .O(N__2422),
            .I(\p.prescaler_1_cry_4 ));
    InMux I__247 (
            .O(N__2419),
            .I(\p.prescaler_1_cry_5 ));
    InMux I__246 (
            .O(N__2416),
            .I(N__2412));
    InMux I__245 (
            .O(N__2415),
            .I(N__2409));
    LocalMux I__244 (
            .O(N__2412),
            .I(\p.prescalerZ0Z_7 ));
    LocalMux I__243 (
            .O(N__2409),
            .I(\p.prescalerZ0Z_7 ));
    InMux I__242 (
            .O(N__2404),
            .I(\p.prescaler_1_cry_6 ));
    InMux I__241 (
            .O(N__2401),
            .I(N__2397));
    InMux I__240 (
            .O(N__2400),
            .I(N__2394));
    LocalMux I__239 (
            .O(N__2397),
            .I(\p.prescalerZ0Z_8 ));
    LocalMux I__238 (
            .O(N__2394),
            .I(\p.prescalerZ0Z_8 ));
    InMux I__237 (
            .O(N__2389),
            .I(\p.prescaler_1_cry_7 ));
    InMux I__236 (
            .O(N__2386),
            .I(N__2382));
    InMux I__235 (
            .O(N__2385),
            .I(N__2379));
    LocalMux I__234 (
            .O(N__2382),
            .I(\p.prescalerZ0Z_9 ));
    LocalMux I__233 (
            .O(N__2379),
            .I(\p.prescalerZ0Z_9 ));
    InMux I__232 (
            .O(N__2374),
            .I(bfn_2_12_0_));
    InMux I__231 (
            .O(N__2371),
            .I(N__2367));
    InMux I__230 (
            .O(N__2370),
            .I(N__2364));
    LocalMux I__229 (
            .O(N__2367),
            .I(\p.prescalerZ0Z_10 ));
    LocalMux I__228 (
            .O(N__2364),
            .I(\p.prescalerZ0Z_10 ));
    InMux I__227 (
            .O(N__2359),
            .I(\p.prescaler_1_cry_9 ));
    InMux I__226 (
            .O(N__2356),
            .I(N__2352));
    InMux I__225 (
            .O(N__2355),
            .I(N__2349));
    LocalMux I__224 (
            .O(N__2352),
            .I(\p.prescalerZ0Z_11 ));
    LocalMux I__223 (
            .O(N__2349),
            .I(\p.prescalerZ0Z_11 ));
    InMux I__222 (
            .O(N__2344),
            .I(\p.prescaler_1_cry_10 ));
    InMux I__221 (
            .O(N__2341),
            .I(N__2338));
    LocalMux I__220 (
            .O(N__2338),
            .I(\p.prescaler12_4_and ));
    InMux I__219 (
            .O(N__2335),
            .I(N__2332));
    LocalMux I__218 (
            .O(N__2332),
            .I(\p.prescaler12_2_and ));
    InMux I__217 (
            .O(N__2329),
            .I(N__2326));
    LocalMux I__216 (
            .O(N__2326),
            .I(\p.prescaler12_6_and ));
    InMux I__215 (
            .O(N__2323),
            .I(N__2320));
    LocalMux I__214 (
            .O(N__2320),
            .I(\p.prescaler12_5_and ));
    InMux I__213 (
            .O(N__2317),
            .I(N__2314));
    LocalMux I__212 (
            .O(N__2314),
            .I(\p.prescaler12_3_and ));
    InMux I__211 (
            .O(N__2311),
            .I(N__2308));
    LocalMux I__210 (
            .O(N__2308),
            .I(N__2305));
    Odrv4 I__209 (
            .O(N__2305),
            .I(\p.prescaler12_1_and ));
    InMux I__208 (
            .O(N__2302),
            .I(N__2297));
    InMux I__207 (
            .O(N__2301),
            .I(N__2292));
    InMux I__206 (
            .O(N__2300),
            .I(N__2292));
    LocalMux I__205 (
            .O(N__2297),
            .I(\p.prescalerZ0Z_2 ));
    LocalMux I__204 (
            .O(N__2292),
            .I(\p.prescalerZ0Z_2 ));
    InMux I__203 (
            .O(N__2287),
            .I(N__2284));
    LocalMux I__202 (
            .O(N__2284),
            .I(\p.prescaler_1_cry_1_THRU_CO ));
    InMux I__201 (
            .O(N__2281),
            .I(\p.prescaler_1_cry_1 ));
    InMux I__200 (
            .O(N__2278),
            .I(\p.prescaler12 ));
    IoInMux I__199 (
            .O(N__2275),
            .I(N__2272));
    LocalMux I__198 (
            .O(N__2272),
            .I(N__2269));
    Odrv12 I__197 (
            .O(N__2269),
            .I(\p.prescaler12_THRU_CO ));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(un1_pulse_len_cry_9),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\p.prescaler_1_cry_8 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\p.prescaler_1_cry_16 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\p.prescaler_1_cry_24 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\p.count_1_cry_8 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\d2.un3_count_cry_8 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\d1.un3_count_cry_8 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\p.CONTROL_PIN_2_cry_9 ),
            .carryinitout(bfn_7_11_0_));
    ICE_GB \p.prescaler12_6_c_RNIPKT  (
            .USERSIGNALTOGLOBALBUFFER(N__2275),
            .GLOBALBUFFEROUTPUT(\p.prescaler12_g ));
    ICE_GB \d2.sync_1_RNIMV5K_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4030),
            .GLOBALBUFFEROUTPUT(\d2.idle_i_g ));
    ICE_GB \d1.sync_1_RNIKI1C_0  (
            .USERSIGNALTOGLOBALBUFFER(N__3499),
            .GLOBALBUFFEROUTPUT(\d1.idle_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \p.prescaler12_0_c_LC_1_11_0 .C_ON=1'b1;
    defparam \p.prescaler12_0_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_0_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_0_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__2584),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\p.prescaler12_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_1_c_LC_1_11_1 .C_ON=1'b1;
    defparam \p.prescaler12_1_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_1_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_1_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__2311),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_0 ),
            .carryout(\p.prescaler12_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_2_c_LC_1_11_2 .C_ON=1'b1;
    defparam \p.prescaler12_2_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_2_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_2_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__2335),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_1 ),
            .carryout(\p.prescaler12_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_3_c_LC_1_11_3 .C_ON=1'b1;
    defparam \p.prescaler12_3_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_3_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_3_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__2317),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_2 ),
            .carryout(\p.prescaler12_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_4_c_LC_1_11_4 .C_ON=1'b1;
    defparam \p.prescaler12_4_c_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_4_c_LC_1_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_4_c_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__2341),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_3 ),
            .carryout(\p.prescaler12_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_5_c_LC_1_11_5 .C_ON=1'b1;
    defparam \p.prescaler12_5_c_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_5_c_LC_1_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_5_c_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__2323),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_4 ),
            .carryout(\p.prescaler12_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_6_c_LC_1_11_6 .C_ON=1'b1;
    defparam \p.prescaler12_6_c_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_6_c_LC_1_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler12_6_c_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__2329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\p.prescaler12_5 ),
            .carryout(\p.prescaler12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_THRU_LUT4_0_LC_1_11_7 .C_ON=1'b0;
    defparam \p.prescaler12_THRU_LUT4_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_THRU_LUT4_0_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \p.prescaler12_THRU_LUT4_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2278),
            .lcout(\p.prescaler12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_4_c_RNO_LC_1_12_0 .C_ON=1'b0;
    defparam \p.prescaler12_4_c_RNO_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_4_c_RNO_LC_1_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.prescaler12_4_c_RNO_LC_1_12_0  (
            .in0(N__2385),
            .in1(N__2355),
            .in2(N__2680),
            .in3(N__2451),
            .lcout(\p.prescaler12_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_2_LC_1_12_1 .C_ON=1'b0;
    defparam \p.prescaler_2_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_2_LC_1_12_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \p.prescaler_2_LC_1_12_1  (
            .in0(N__2287),
            .in1(N__2301),
            .in2(_gnd_net_),
            .in3(N__4439),
            .lcout(\p.prescalerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4812),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_2_c_RNO_LC_1_12_3 .C_ON=1'b0;
    defparam \p.prescaler12_2_c_RNO_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_2_c_RNO_LC_1_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.prescaler12_2_c_RNO_LC_1_12_3  (
            .in0(N__2499),
            .in1(N__2559),
            .in2(N__2623),
            .in3(N__2574),
            .lcout(\p.prescaler12_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_6_c_RNO_LC_1_12_4 .C_ON=1'b0;
    defparam \p.prescaler12_6_c_RNO_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_6_c_RNO_LC_1_12_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \p.prescaler12_6_c_RNO_LC_1_12_4  (
            .in0(N__2466),
            .in1(N__2514),
            .in2(_gnd_net_),
            .in3(N__2415),
            .lcout(\p.prescaler12_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_5_c_RNO_LC_1_12_6 .C_ON=1'b0;
    defparam \p.prescaler12_5_c_RNO_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_5_c_RNO_LC_1_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.prescaler12_5_c_RNO_LC_1_12_6  (
            .in0(N__2529),
            .in1(N__2400),
            .in2(N__2644),
            .in3(N__2436),
            .lcout(\p.prescaler12_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_3_c_RNO_LC_1_12_7 .C_ON=1'b0;
    defparam \p.prescaler12_3_c_RNO_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_3_c_RNO_LC_1_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.prescaler12_3_c_RNO_LC_1_12_7  (
            .in0(N__2370),
            .in1(N__2485),
            .in2(N__2662),
            .in3(N__2300),
            .lcout(\p.prescaler12_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_1_c_RNO_LC_1_13_1 .C_ON=1'b0;
    defparam \p.prescaler12_1_c_RNO_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_1_c_RNO_LC_1_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.prescaler12_1_c_RNO_LC_1_13_1  (
            .in0(N__2694),
            .in1(N__2709),
            .in2(N__2599),
            .in3(N__2544),
            .lcout(\p.prescaler12_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_1_cry_1_c_LC_2_11_0 .C_ON=1'b1;
    defparam \p.prescaler_1_cry_1_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \p.prescaler_1_cry_1_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.prescaler_1_cry_1_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__2761),
            .in2(N__2743),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\p.prescaler_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_1_cry_1_THRU_LUT4_0_LC_2_11_1 .C_ON=1'b1;
    defparam \p.prescaler_1_cry_1_THRU_LUT4_0_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \p.prescaler_1_cry_1_THRU_LUT4_0_LC_2_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \p.prescaler_1_cry_1_THRU_LUT4_0_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__2302),
            .in2(_gnd_net_),
            .in3(N__2281),
            .lcout(\p.prescaler_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_1 ),
            .carryout(\p.prescaler_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_3_LC_2_11_2 .C_ON=1'b1;
    defparam \p.prescaler_3_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_3_LC_2_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_3_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__2452),
            .in2(_gnd_net_),
            .in3(N__2440),
            .lcout(\p.prescalerZ0Z_3 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_2 ),
            .carryout(\p.prescaler_1_cry_3 ),
            .clk(N__4813),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_4_LC_2_11_3 .C_ON=1'b1;
    defparam \p.prescaler_4_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_4_LC_2_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_4_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__2437),
            .in2(_gnd_net_),
            .in3(N__2425),
            .lcout(\p.prescalerZ0Z_4 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_3 ),
            .carryout(\p.prescaler_1_cry_4 ),
            .clk(N__4813),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_1_cry_4_THRU_LUT4_0_LC_2_11_4 .C_ON=1'b1;
    defparam \p.prescaler_1_cry_4_THRU_LUT4_0_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \p.prescaler_1_cry_4_THRU_LUT4_0_LC_2_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \p.prescaler_1_cry_4_THRU_LUT4_0_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__2776),
            .in2(_gnd_net_),
            .in3(N__2422),
            .lcout(\p.prescaler_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_4 ),
            .carryout(\p.prescaler_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_1_cry_5_THRU_LUT4_0_LC_2_11_5 .C_ON=1'b1;
    defparam \p.prescaler_1_cry_5_THRU_LUT4_0_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \p.prescaler_1_cry_5_THRU_LUT4_0_LC_2_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \p.prescaler_1_cry_5_THRU_LUT4_0_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__2801),
            .in2(_gnd_net_),
            .in3(N__2419),
            .lcout(\p.prescaler_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_5 ),
            .carryout(\p.prescaler_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_7_LC_2_11_6 .C_ON=1'b1;
    defparam \p.prescaler_7_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_7_LC_2_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_7_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__2416),
            .in2(_gnd_net_),
            .in3(N__2404),
            .lcout(\p.prescalerZ0Z_7 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_6 ),
            .carryout(\p.prescaler_1_cry_7 ),
            .clk(N__4813),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_8_LC_2_11_7 .C_ON=1'b1;
    defparam \p.prescaler_8_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_8_LC_2_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__2401),
            .in2(_gnd_net_),
            .in3(N__2389),
            .lcout(\p.prescalerZ0Z_8 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_7 ),
            .carryout(\p.prescaler_1_cry_8 ),
            .clk(N__4813),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_9_LC_2_12_0 .C_ON=1'b1;
    defparam \p.prescaler_9_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_9_LC_2_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_9_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__2386),
            .in2(_gnd_net_),
            .in3(N__2374),
            .lcout(\p.prescalerZ0Z_9 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\p.prescaler_1_cry_9 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_10_LC_2_12_1 .C_ON=1'b1;
    defparam \p.prescaler_10_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_10_LC_2_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_10_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__2371),
            .in2(_gnd_net_),
            .in3(N__2359),
            .lcout(\p.prescalerZ0Z_10 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_9 ),
            .carryout(\p.prescaler_1_cry_10 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_11_LC_2_12_2 .C_ON=1'b1;
    defparam \p.prescaler_11_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_11_LC_2_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_11_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__2356),
            .in2(_gnd_net_),
            .in3(N__2344),
            .lcout(\p.prescalerZ0Z_11 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_10 ),
            .carryout(\p.prescaler_1_cry_11 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_12_LC_2_12_3 .C_ON=1'b1;
    defparam \p.prescaler_12_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_12_LC_2_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_12_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__2575),
            .in2(_gnd_net_),
            .in3(N__2563),
            .lcout(\p.prescalerZ0Z_12 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_11 ),
            .carryout(\p.prescaler_1_cry_12 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_13_LC_2_12_4 .C_ON=1'b1;
    defparam \p.prescaler_13_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_13_LC_2_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_13_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__2560),
            .in2(_gnd_net_),
            .in3(N__2548),
            .lcout(\p.prescalerZ0Z_13 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_12 ),
            .carryout(\p.prescaler_1_cry_13 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_14_LC_2_12_5 .C_ON=1'b1;
    defparam \p.prescaler_14_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_14_LC_2_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_14_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__2545),
            .in2(_gnd_net_),
            .in3(N__2533),
            .lcout(\p.prescalerZ0Z_14 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_13 ),
            .carryout(\p.prescaler_1_cry_14 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_15_LC_2_12_6 .C_ON=1'b1;
    defparam \p.prescaler_15_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_15_LC_2_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_15_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__2530),
            .in2(_gnd_net_),
            .in3(N__2518),
            .lcout(\p.prescalerZ0Z_15 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_14 ),
            .carryout(\p.prescaler_1_cry_15 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_16_LC_2_12_7 .C_ON=1'b1;
    defparam \p.prescaler_16_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_16_LC_2_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_16_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__2515),
            .in2(_gnd_net_),
            .in3(N__2503),
            .lcout(\p.prescalerZ0Z_16 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_15 ),
            .carryout(\p.prescaler_1_cry_16 ),
            .clk(N__4809),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_17_LC_2_13_0 .C_ON=1'b1;
    defparam \p.prescaler_17_LC_2_13_0 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_17_LC_2_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_17_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__2500),
            .in2(_gnd_net_),
            .in3(N__2488),
            .lcout(\p.prescalerZ0Z_17 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\p.prescaler_1_cry_17 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_18_LC_2_13_1 .C_ON=1'b1;
    defparam \p.prescaler_18_LC_2_13_1 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_18_LC_2_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_18_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__2484),
            .in2(_gnd_net_),
            .in3(N__2470),
            .lcout(\p.prescalerZ0Z_18 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_17 ),
            .carryout(\p.prescaler_1_cry_18 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_19_LC_2_13_2 .C_ON=1'b1;
    defparam \p.prescaler_19_LC_2_13_2 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_19_LC_2_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_19_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__2467),
            .in2(_gnd_net_),
            .in3(N__2455),
            .lcout(\p.prescalerZ0Z_19 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_18 ),
            .carryout(\p.prescaler_1_cry_19 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_20_LC_2_13_3 .C_ON=1'b1;
    defparam \p.prescaler_20_LC_2_13_3 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_20_LC_2_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_20_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__2710),
            .in2(_gnd_net_),
            .in3(N__2698),
            .lcout(\p.prescalerZ0Z_20 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_19 ),
            .carryout(\p.prescaler_1_cry_20 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_21_LC_2_13_4 .C_ON=1'b1;
    defparam \p.prescaler_21_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_21_LC_2_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_21_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__2695),
            .in2(_gnd_net_),
            .in3(N__2683),
            .lcout(\p.prescalerZ0Z_21 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_20 ),
            .carryout(\p.prescaler_1_cry_21 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_22_LC_2_13_5 .C_ON=1'b1;
    defparam \p.prescaler_22_LC_2_13_5 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_22_LC_2_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_22_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__2679),
            .in2(_gnd_net_),
            .in3(N__2665),
            .lcout(\p.prescalerZ0Z_22 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_21 ),
            .carryout(\p.prescaler_1_cry_22 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_23_LC_2_13_6 .C_ON=1'b1;
    defparam \p.prescaler_23_LC_2_13_6 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_23_LC_2_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_23_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__2661),
            .in2(_gnd_net_),
            .in3(N__2647),
            .lcout(\p.prescalerZ0Z_23 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_22 ),
            .carryout(\p.prescaler_1_cry_23 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_24_LC_2_13_7 .C_ON=1'b1;
    defparam \p.prescaler_24_LC_2_13_7 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_24_LC_2_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_24_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__2640),
            .in2(_gnd_net_),
            .in3(N__2626),
            .lcout(\p.prescalerZ0Z_24 ),
            .ltout(),
            .carryin(\p.prescaler_1_cry_23 ),
            .carryout(\p.prescaler_1_cry_24 ),
            .clk(N__4808),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_25_LC_2_14_0 .C_ON=1'b1;
    defparam \p.prescaler_25_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_25_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.prescaler_25_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__2619),
            .in2(_gnd_net_),
            .in3(N__2605),
            .lcout(\p.prescalerZ0Z_25 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\p.prescaler_1_cry_25 ),
            .clk(N__4805),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_26_LC_2_14_1 .C_ON=1'b0;
    defparam \p.prescaler_26_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_26_LC_2_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \p.prescaler_26_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__2598),
            .in2(_gnd_net_),
            .in3(N__2602),
            .lcout(\p.prescalerZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4805),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_0_LC_3_11_2 .C_ON=1'b0;
    defparam \p.prescaler_0_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_0_LC_3_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \p.prescaler_0_LC_3_11_2  (
            .in0(N__2759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\p.prescalerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler12_0_c_RNO_LC_3_11_3 .C_ON=1'b0;
    defparam \p.prescaler12_0_c_RNO_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \p.prescaler12_0_c_RNO_LC_3_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \p.prescaler12_0_c_RNO_LC_3_11_3  (
            .in0(N__2774),
            .in1(N__2738),
            .in2(N__2802),
            .in3(N__2758),
            .lcout(\p.prescaler12_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_6_LC_3_11_5 .C_ON=1'b0;
    defparam \p.prescaler_6_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_6_LC_3_11_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \p.prescaler_6_LC_3_11_5  (
            .in0(N__4441),
            .in1(_gnd_net_),
            .in2(N__2803),
            .in3(N__2809),
            .lcout(\p.prescalerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_5_LC_3_11_6 .C_ON=1'b0;
    defparam \p.prescaler_5_LC_3_11_6 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_5_LC_3_11_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \p.prescaler_5_LC_3_11_6  (
            .in0(N__2782),
            .in1(N__2775),
            .in2(_gnd_net_),
            .in3(N__4440),
            .lcout(\p.prescalerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.prescaler_1_LC_3_11_7 .C_ON=1'b0;
    defparam \p.prescaler_1_LC_3_11_7 .SEQ_MODE=4'b1000;
    defparam \p.prescaler_1_LC_3_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \p.prescaler_1_LC_3_11_7  (
            .in0(_gnd_net_),
            .in1(N__2739),
            .in2(_gnd_net_),
            .in3(N__2760),
            .lcout(\p.prescalerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4810),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_6_LC_7_7_5 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_6_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_6_LC_7_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \d2.state_RNIPC4P3_6_LC_7_7_5  (
            .in0(N__3456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4084),
            .lcout(state_RNIPC4P3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_LC_7_7_6 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_LC_7_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__4076),
            .in2(_gnd_net_),
            .in3(N__3455),
            .lcout(state_RNIPC4P3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_pulse_len_cry_2_c_LC_7_8_0.C_ON=1'b1;
    defparam un1_pulse_len_cry_2_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam un1_pulse_len_cry_2_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_pulse_len_cry_2_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__3331),
            .in2(N__3307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(un1_pulse_len_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_3_LC_7_8_1.C_ON=1'b1;
    defparam pulse_len_3_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam pulse_len_3_LC_7_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_3_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__2725),
            .in2(N__2946),
            .in3(N__2719),
            .lcout(pulse_lenZ0Z_3),
            .ltout(),
            .carryin(un1_pulse_len_cry_2),
            .carryout(un1_pulse_len_cry_3),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_4_LC_7_8_2.C_ON=1'b1;
    defparam pulse_len_4_LC_7_8_2.SEQ_MODE=4'b1000;
    defparam pulse_len_4_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_4_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__3361),
            .in2(N__2919),
            .in3(N__2716),
            .lcout(pulse_lenZ0Z_4),
            .ltout(),
            .carryin(un1_pulse_len_cry_3),
            .carryout(un1_pulse_len_cry_4),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_5_LC_7_8_3.C_ON=1'b1;
    defparam pulse_len_5_LC_7_8_3.SEQ_MODE=4'b1000;
    defparam pulse_len_5_LC_7_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_5_LC_7_8_3 (
            .in0(_gnd_net_),
            .in1(N__2886),
            .in2(N__3370),
            .in3(N__2713),
            .lcout(pulse_lenZ0Z_5),
            .ltout(),
            .carryin(un1_pulse_len_cry_4),
            .carryout(un1_pulse_len_cry_5),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_6_LC_7_8_4.C_ON=1'b1;
    defparam pulse_len_6_LC_7_8_4.SEQ_MODE=4'b1000;
    defparam pulse_len_6_LC_7_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_6_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__2862),
            .in2(N__3487),
            .in3(N__2842),
            .lcout(pulse_lenZ0Z_6),
            .ltout(),
            .carryin(un1_pulse_len_cry_5),
            .carryout(un1_pulse_len_cry_6),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_7_LC_7_8_5.C_ON=1'b1;
    defparam pulse_len_7_LC_7_8_5.SEQ_MODE=4'b1000;
    defparam pulse_len_7_LC_7_8_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_7_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(N__3298),
            .in2(N__3192),
            .in3(N__2839),
            .lcout(pulse_lenZ0Z_7),
            .ltout(),
            .carryin(un1_pulse_len_cry_6),
            .carryout(un1_pulse_len_cry_7),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_8_LC_7_8_6.C_ON=1'b1;
    defparam pulse_len_8_LC_7_8_6.SEQ_MODE=4'b1000;
    defparam pulse_len_8_LC_7_8_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_8_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(N__2836),
            .in2(N__3165),
            .in3(N__2830),
            .lcout(pulse_lenZ0Z_8),
            .ltout(),
            .carryin(un1_pulse_len_cry_7),
            .carryout(un1_pulse_len_cry_8),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_9_LC_7_8_7.C_ON=1'b1;
    defparam pulse_len_9_LC_7_8_7.SEQ_MODE=4'b1000;
    defparam pulse_len_9_LC_7_8_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_9_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(N__3355),
            .in2(N__3136),
            .in3(N__2827),
            .lcout(pulse_lenZ0Z_9),
            .ltout(),
            .carryin(un1_pulse_len_cry_8),
            .carryout(un1_pulse_len_cry_9),
            .clk(N__4806),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_10_LC_7_9_0.C_ON=1'b1;
    defparam pulse_len_10_LC_7_9_0.SEQ_MODE=4'b1000;
    defparam pulse_len_10_LC_7_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_10_LC_7_9_0 (
            .in0(_gnd_net_),
            .in1(N__3478),
            .in2(N__3108),
            .in3(N__2824),
            .lcout(pulse_lenZ0Z_10),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(un1_pulse_len_cry_10),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_11_LC_7_9_1.C_ON=1'b1;
    defparam pulse_len_11_LC_7_9_1.SEQ_MODE=4'b1000;
    defparam pulse_len_11_LC_7_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_11_LC_7_9_1 (
            .in0(_gnd_net_),
            .in1(N__3415),
            .in2(N__3078),
            .in3(N__2821),
            .lcout(pulse_lenZ0Z_11),
            .ltout(),
            .carryin(un1_pulse_len_cry_10),
            .carryout(un1_pulse_len_cry_11),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_12_LC_7_9_2.C_ON=1'b1;
    defparam pulse_len_12_LC_7_9_2.SEQ_MODE=4'b1000;
    defparam pulse_len_12_LC_7_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_12_LC_7_9_2 (
            .in0(_gnd_net_),
            .in1(N__2962),
            .in2(N__3051),
            .in3(N__2818),
            .lcout(pulse_lenZ0Z_12),
            .ltout(),
            .carryin(un1_pulse_len_cry_11),
            .carryout(un1_pulse_len_cry_12),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_13_LC_7_9_3.C_ON=1'b1;
    defparam pulse_len_13_LC_7_9_3.SEQ_MODE=4'b1000;
    defparam pulse_len_13_LC_7_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_13_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(N__2968),
            .in2(N__3024),
            .in3(N__2815),
            .lcout(pulse_lenZ0Z_13),
            .ltout(),
            .carryin(un1_pulse_len_cry_12),
            .carryout(un1_pulse_len_cry_13),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_14_LC_7_9_4.C_ON=1'b1;
    defparam pulse_len_14_LC_7_9_4.SEQ_MODE=4'b1000;
    defparam pulse_len_14_LC_7_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 pulse_len_14_LC_7_9_4 (
            .in0(_gnd_net_),
            .in1(N__3472),
            .in2(N__2997),
            .in3(N__2812),
            .lcout(pulse_lenZ0Z_14),
            .ltout(),
            .carryin(un1_pulse_len_cry_13),
            .carryout(un1_pulse_len_cry_14),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_15_LC_7_9_5.C_ON=1'b0;
    defparam pulse_len_15_LC_7_9_5.SEQ_MODE=4'b1000;
    defparam pulse_len_15_LC_7_9_5.LUT_INIT=16'b1000011101111000;
    LogicCell40 pulse_len_15_LC_7_9_5 (
            .in0(N__4117),
            .in1(N__3466),
            .in2(N__3264),
            .in3(N__2971),
            .lcout(pulse_lenZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4802),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_4_LC_7_9_6 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_4_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_4_LC_7_9_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \d2.state_RNIPC4P3_4_LC_7_9_6  (
            .in0(N__3465),
            .in1(_gnd_net_),
            .in2(N__4116),
            .in3(_gnd_net_),
            .lcout(state_RNIPC4P3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_7_LC_7_9_7 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_7_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_7_LC_7_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_7_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__4108),
            .in2(_gnd_net_),
            .in3(N__3464),
            .lcout(state_RNIPC4P3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_2_c_inv_LC_7_10_0 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_2_c_inv_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_2_c_inv_LC_7_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_2_c_inv_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__2956),
            .in2(N__3340),
            .in3(N__3622),
            .lcout(\p.count_i_2 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\p.CONTROL_PIN_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_3_c_inv_LC_7_10_1 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_3_c_inv_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_3_c_inv_LC_7_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_3_c_inv_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__2926),
            .in2(N__2950),
            .in3(N__3643),
            .lcout(\p.count_i_3 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_2 ),
            .carryout(\p.CONTROL_PIN_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_4_c_inv_LC_7_10_2 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_4_c_inv_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_4_c_inv_LC_7_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_4_c_inv_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__2899),
            .in2(N__2920),
            .in3(N__3703),
            .lcout(\p.count_i_4 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_3 ),
            .carryout(\p.CONTROL_PIN_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_5_c_inv_LC_7_10_3 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_5_c_inv_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_5_c_inv_LC_7_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_5_c_inv_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__2872),
            .in2(N__2893),
            .in3(N__3790),
            .lcout(\p.count_i_5 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_4 ),
            .carryout(\p.CONTROL_PIN_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_6_c_inv_LC_7_10_4 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_6_c_inv_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_6_c_inv_LC_7_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_6_c_inv_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__2848),
            .in2(N__2866),
            .in3(N__3877),
            .lcout(\p.count_i_6 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_5 ),
            .carryout(\p.CONTROL_PIN_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_7_c_inv_LC_7_10_5 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_7_c_inv_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_7_c_inv_LC_7_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \p.CONTROL_PIN_2_cry_7_c_inv_LC_7_10_5  (
            .in0(N__3835),
            .in1(N__3172),
            .in2(N__3196),
            .in3(_gnd_net_),
            .lcout(\p.count_i_7 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_6 ),
            .carryout(\p.CONTROL_PIN_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_8_c_inv_LC_7_10_6 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_8_c_inv_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_8_c_inv_LC_7_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_8_c_inv_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__3142),
            .in2(N__3166),
            .in3(N__3922),
            .lcout(\p.count_i_8 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_7 ),
            .carryout(\p.CONTROL_PIN_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_9_c_inv_LC_7_10_7 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_9_c_inv_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_9_c_inv_LC_7_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_9_c_inv_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__3135),
            .in2(N__3118),
            .in3(N__3748),
            .lcout(\p.count_i_9 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_8 ),
            .carryout(\p.CONTROL_PIN_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_10_c_inv_LC_7_11_0 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_10_c_inv_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_10_c_inv_LC_7_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_10_c_inv_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__3088),
            .in2(N__3109),
            .in3(N__3769),
            .lcout(\p.count_i_10 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\p.CONTROL_PIN_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_11_c_inv_LC_7_11_1 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_11_c_inv_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_11_c_inv_LC_7_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_11_c_inv_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__3058),
            .in2(N__3082),
            .in3(N__3726),
            .lcout(\p.count_i_11 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_10 ),
            .carryout(\p.CONTROL_PIN_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_12_c_inv_LC_7_11_2 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_12_c_inv_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_12_c_inv_LC_7_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_12_c_inv_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__3031),
            .in2(N__3052),
            .in3(N__3856),
            .lcout(\p.count_i_12 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_11 ),
            .carryout(\p.CONTROL_PIN_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_13_c_inv_LC_7_11_3 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_13_c_inv_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_13_c_inv_LC_7_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_13_c_inv_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__3004),
            .in2(N__3025),
            .in3(N__3813),
            .lcout(\p.count_i_13 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_12 ),
            .carryout(\p.CONTROL_PIN_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_14_c_inv_LC_7_11_4 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_14_c_inv_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_14_c_inv_LC_7_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.CONTROL_PIN_2_cry_14_c_inv_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__2977),
            .in2(N__2998),
            .in3(N__3943),
            .lcout(\p.count_i_14 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_13 ),
            .carryout(\p.CONTROL_PIN_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_2_cry_15_c_inv_LC_7_11_5 .C_ON=1'b1;
    defparam \p.CONTROL_PIN_2_cry_15_c_inv_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \p.CONTROL_PIN_2_cry_15_c_inv_LC_7_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \p.CONTROL_PIN_2_cry_15_c_inv_LC_7_11_5  (
            .in0(N__3901),
            .in1(N__3244),
            .in2(N__3268),
            .in3(_gnd_net_),
            .lcout(\p.count_i_15 ),
            .ltout(),
            .carryin(\p.CONTROL_PIN_2_cry_14 ),
            .carryout(\p.CONTROL_PIN_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.CONTROL_PIN_LC_7_11_6 .C_ON=1'b0;
    defparam \p.CONTROL_PIN_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \p.CONTROL_PIN_LC_7_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \p.CONTROL_PIN_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3238),
            .lcout(CONTROL_PIN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4797),
            .ce(N__4427),
            .sr(_gnd_net_));
    defparam \p.count_1_cry_1_c_LC_7_12_0 .C_ON=1'b1;
    defparam \p.count_1_cry_1_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \p.count_1_cry_1_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \p.count_1_cry_1_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__4465),
            .in2(N__4492),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\p.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.count_2_LC_7_12_1 .C_ON=1'b1;
    defparam \p.count_2_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \p.count_2_LC_7_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_2_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__3621),
            .in2(_gnd_net_),
            .in3(N__3214),
            .lcout(\p.countZ0Z_2 ),
            .ltout(),
            .carryin(\p.count_1_cry_1 ),
            .carryout(\p.count_1_cry_2 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_3_LC_7_12_2 .C_ON=1'b1;
    defparam \p.count_3_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \p.count_3_LC_7_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_3_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__3642),
            .in2(_gnd_net_),
            .in3(N__3211),
            .lcout(\p.countZ0Z_3 ),
            .ltout(),
            .carryin(\p.count_1_cry_2 ),
            .carryout(\p.count_1_cry_3 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_4_LC_7_12_3 .C_ON=1'b1;
    defparam \p.count_4_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \p.count_4_LC_7_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_4_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__3702),
            .in2(_gnd_net_),
            .in3(N__3208),
            .lcout(\p.countZ0Z_4 ),
            .ltout(),
            .carryin(\p.count_1_cry_3 ),
            .carryout(\p.count_1_cry_4 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_5_LC_7_12_4 .C_ON=1'b1;
    defparam \p.count_5_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \p.count_5_LC_7_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \p.count_5_LC_7_12_4  (
            .in0(N__3665),
            .in1(N__3789),
            .in2(_gnd_net_),
            .in3(N__3205),
            .lcout(\p.countZ0Z_5 ),
            .ltout(),
            .carryin(\p.count_1_cry_4 ),
            .carryout(\p.count_1_cry_5 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_6_LC_7_12_5 .C_ON=1'b1;
    defparam \p.count_6_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \p.count_6_LC_7_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_6_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__3876),
            .in2(_gnd_net_),
            .in3(N__3202),
            .lcout(\p.countZ0Z_6 ),
            .ltout(),
            .carryin(\p.count_1_cry_5 ),
            .carryout(\p.count_1_cry_6 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_7_LC_7_12_6 .C_ON=1'b1;
    defparam \p.count_7_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \p.count_7_LC_7_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_7_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__3834),
            .in2(_gnd_net_),
            .in3(N__3199),
            .lcout(\p.countZ0Z_7 ),
            .ltout(),
            .carryin(\p.count_1_cry_6 ),
            .carryout(\p.count_1_cry_7 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_8_LC_7_12_7 .C_ON=1'b1;
    defparam \p.count_8_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \p.count_8_LC_7_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_8_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__3921),
            .in2(_gnd_net_),
            .in3(N__3292),
            .lcout(\p.countZ0Z_8 ),
            .ltout(),
            .carryin(\p.count_1_cry_7 ),
            .carryout(\p.count_1_cry_8 ),
            .clk(N__4793),
            .ce(N__4428),
            .sr(_gnd_net_));
    defparam \p.count_9_LC_7_13_0 .C_ON=1'b1;
    defparam \p.count_9_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \p.count_9_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \p.count_9_LC_7_13_0  (
            .in0(N__3664),
            .in1(N__3747),
            .in2(_gnd_net_),
            .in3(N__3289),
            .lcout(\p.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\p.count_1_cry_9 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_10_LC_7_13_1 .C_ON=1'b1;
    defparam \p.count_10_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \p.count_10_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \p.count_10_LC_7_13_1  (
            .in0(N__3666),
            .in1(N__3768),
            .in2(_gnd_net_),
            .in3(N__3286),
            .lcout(\p.countZ0Z_10 ),
            .ltout(),
            .carryin(\p.count_1_cry_9 ),
            .carryout(\p.count_1_cry_10 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_11_LC_7_13_2 .C_ON=1'b1;
    defparam \p.count_11_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \p.count_11_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \p.count_11_LC_7_13_2  (
            .in0(N__3663),
            .in1(N__3725),
            .in2(_gnd_net_),
            .in3(N__3283),
            .lcout(\p.countZ0Z_11 ),
            .ltout(),
            .carryin(\p.count_1_cry_10 ),
            .carryout(\p.count_1_cry_11 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_12_LC_7_13_3 .C_ON=1'b1;
    defparam \p.count_12_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \p.count_12_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_12_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__3855),
            .in2(_gnd_net_),
            .in3(N__3280),
            .lcout(\p.countZ0Z_12 ),
            .ltout(),
            .carryin(\p.count_1_cry_11 ),
            .carryout(\p.count_1_cry_12 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_13_LC_7_13_4 .C_ON=1'b1;
    defparam \p.count_13_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \p.count_13_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \p.count_13_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__3812),
            .in2(_gnd_net_),
            .in3(N__3277),
            .lcout(\p.countZ0Z_13 ),
            .ltout(),
            .carryin(\p.count_1_cry_12 ),
            .carryout(\p.count_1_cry_13 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_14_LC_7_13_5 .C_ON=1'b1;
    defparam \p.count_14_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \p.count_14_LC_7_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \p.count_14_LC_7_13_5  (
            .in0(N__3667),
            .in1(N__3942),
            .in2(_gnd_net_),
            .in3(N__3274),
            .lcout(\p.countZ0Z_14 ),
            .ltout(),
            .carryin(\p.count_1_cry_13 ),
            .carryout(\p.count_1_cry_14 ),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \p.count_15_LC_7_13_6 .C_ON=1'b0;
    defparam \p.count_15_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \p.count_15_LC_7_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \p.count_15_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__3899),
            .in2(_gnd_net_),
            .in3(N__3271),
            .lcout(\p.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4792),
            .ce(N__4429),
            .sr(_gnd_net_));
    defparam \d2.state_LC_8_7_0 .C_ON=1'b0;
    defparam \d2.state_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \d2.state_LC_8_7_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \d2.state_LC_8_7_0  (
            .in0(N__3459),
            .in1(_gnd_net_),
            .in2(N__4102),
            .in3(_gnd_net_),
            .lcout(d2_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4807),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_0_LC_8_7_3 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_0_LC_8_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_0_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__4077),
            .in2(_gnd_net_),
            .in3(N__3457),
            .lcout(state_RNIPC4P3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_2_LC_8_7_4 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_2_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_2_LC_8_7_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \d2.state_RNIPC4P3_2_LC_8_7_4  (
            .in0(N__3458),
            .in1(_gnd_net_),
            .in2(N__4101),
            .in3(_gnd_net_),
            .lcout(state_RNIPC4P3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pulse_len_2_LC_8_8_0.C_ON=1'b0;
    defparam pulse_len_2_LC_8_8_0.SEQ_MODE=4'b1000;
    defparam pulse_len_2_LC_8_8_0.LUT_INIT=16'b0000101011110101;
    LogicCell40 pulse_len_2_LC_8_8_0 (
            .in0(N__3385),
            .in1(_gnd_net_),
            .in2(N__3403),
            .in3(N__3335),
            .lcout(pulse_lenZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4803),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNINDU8_0_LC_8_8_1 .C_ON=1'b0;
    defparam \d2.count_RNINDU8_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNINDU8_0_LC_8_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \d2.count_RNINDU8_0_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__4396),
            .in2(_gnd_net_),
            .in3(N__4174),
            .lcout(),
            .ltout(\d2.trans_up_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_RNI3PR51_LC_8_8_2 .C_ON=1'b0;
    defparam \d2.sync_1_RNI3PR51_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \d2.sync_1_RNI3PR51_LC_8_8_2 .LUT_INIT=16'b1011111101111111;
    LogicCell40 \d2.sync_1_RNI3PR51_LC_8_8_2  (
            .in0(N__4128),
            .in1(N__4370),
            .in2(N__3349),
            .in3(N__4073),
            .lcout(),
            .ltout(\d2.trans_up_1_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIK9TB3_10_LC_8_8_3 .C_ON=1'b0;
    defparam \d2.count_RNIK9TB3_10_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIK9TB3_10_LC_8_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \d2.count_RNIK9TB3_10_LC_8_8_3  (
            .in0(N__3595),
            .in1(N__3583),
            .in2(N__3346),
            .in3(N__4186),
            .lcout(d2_trans_up_1),
            .ltout(d2_trans_up_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_9_LC_8_8_4 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_9_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_9_LC_8_8_4 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \d2.state_RNIPC4P3_9_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3343),
            .in3(N__4074),
            .lcout(s_dn_i),
            .ltout(s_dn_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_pulse_len_cry_2_c_RNO_LC_8_8_5.C_ON=1'b0;
    defparam un1_pulse_len_cry_2_c_RNO_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam un1_pulse_len_cry_2_c_RNO_LC_8_8_5.LUT_INIT=16'b1111111100001111;
    LogicCell40 un1_pulse_len_cry_2_c_RNO_LC_8_8_5 (
            .in0(N__3336),
            .in1(_gnd_net_),
            .in2(N__3310),
            .in3(N__3398),
            .lcout(un1_pulse_len_cry_2_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_3_LC_8_8_6 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_3_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_3_LC_8_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_3_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__4075),
            .in2(_gnd_net_),
            .in3(N__3460),
            .lcout(state_RNIPC4P3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIU5D07_LC_8_8_7 .C_ON=1'b0;
    defparam \d2.state_RNIU5D07_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIU5D07_LC_8_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIU5D07_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__3399),
            .in2(_gnd_net_),
            .in3(N__3384),
            .lcout(state_RNIU5D07),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_1_LC_8_9_0 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_1_LC_8_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_1_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__4103),
            .in2(_gnd_net_),
            .in3(N__3461),
            .lcout(state_RNIPC4P3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_8_LC_8_9_1 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_8_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_8_LC_8_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \d2.state_RNIPC4P3_8_LC_8_9_1  (
            .in0(N__3463),
            .in1(_gnd_net_),
            .in2(N__4115),
            .in3(_gnd_net_),
            .lcout(state_RNIPC4P3_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIPC4P3_5_LC_8_9_2 .C_ON=1'b0;
    defparam \d2.state_RNIPC4P3_5_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIPC4P3_5_LC_8_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \d2.state_RNIPC4P3_5_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__4104),
            .in2(_gnd_net_),
            .in3(N__3462),
            .lcout(state_RNIPC4P3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_LC_8_9_3 .C_ON=1'b0;
    defparam \d1.sync_1_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \d1.sync_1_LC_8_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d1.sync_1_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4822),
            .lcout(\d1.syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4800),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI2PCE_3_LC_8_9_4 .C_ON=1'b0;
    defparam \d1.count_RNI2PCE_3_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI2PCE_3_LC_8_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI2PCE_3_LC_8_9_4  (
            .in0(N__4323),
            .in1(N__4338),
            .in2(N__4309),
            .in3(N__4353),
            .lcout(),
            .ltout(\d1.count_RNI2PCEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI23S21_3_LC_8_9_5 .C_ON=1'b0;
    defparam \d1.count_RNI23S21_3_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI23S21_3_LC_8_9_5 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \d1.count_RNI23S21_3_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__3571),
            .in2(N__3409),
            .in3(_gnd_net_),
            .lcout(\d1.trans_up_1_14 ),
            .ltout(\d1.trans_up_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI5P873_7_LC_8_9_6 .C_ON=1'b0;
    defparam \d1.count_RNI5P873_7_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI5P873_7_LC_8_9_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \d1.count_RNI5P873_7_LC_8_9_6  (
            .in0(N__3535),
            .in1(N__3552),
            .in2(N__3406),
            .in3(N__3541),
            .lcout(s_up),
            .ltout(s_up_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNIU5D07_0_LC_8_9_7 .C_ON=1'b0;
    defparam \d2.state_RNIU5D07_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNIU5D07_0_LC_8_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \d2.state_RNIU5D07_0_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3388),
            .in3(N__3383),
            .lcout(state_RNIU5D07_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI0AFK_16_LC_8_10_0 .C_ON=1'b0;
    defparam \d1.count_RNI0AFK_16_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI0AFK_16_LC_8_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI0AFK_16_LC_8_10_0  (
            .in0(N__3957),
            .in1(N__4004),
            .in2(N__4522),
            .in3(N__4539),
            .lcout(\d1.trans_up_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_RNI5IAP_LC_8_10_1 .C_ON=1'b0;
    defparam \d1.sync_1_RNI5IAP_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \d1.sync_1_RNI5IAP_LC_8_10_1 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \d1.sync_1_RNI5IAP_LC_8_10_1  (
            .in0(N__3526),
            .in1(N__4554),
            .in2(N__3514),
            .in3(N__4569),
            .lcout(\d1.trans_up_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNO_1_LC_8_10_2 .C_ON=1'b0;
    defparam \d1.state_RNO_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNO_1_LC_8_10_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.state_RNO_1_LC_8_10_2  (
            .in0(N__4290),
            .in1(N__4251),
            .in2(N__4233),
            .in3(N__4272),
            .lcout(),
            .ltout(\d1.trans_up_1_13_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNO_0_LC_8_10_3 .C_ON=1'b0;
    defparam \d1.state_RNO_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNO_0_LC_8_10_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \d1.state_RNO_0_LC_8_10_3  (
            .in0(N__3979),
            .in1(N__4589),
            .in2(N__3565),
            .in3(N__4203),
            .lcout(),
            .ltout(\d1.trans_up_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_LC_8_10_4 .C_ON=1'b0;
    defparam \d1.state_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \d1.state_LC_8_10_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \d1.state_LC_8_10_4  (
            .in0(N__3562),
            .in1(N__3529),
            .in2(N__3556),
            .in3(N__3553),
            .lcout(\d1.stateZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4798),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIP9EH_7_LC_8_10_5 .C_ON=1'b0;
    defparam \d1.count_RNIP9EH_7_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIP9EH_7_LC_8_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNIP9EH_7_LC_8_10_5  (
            .in0(N__4250),
            .in1(N__4271),
            .in2(N__4234),
            .in3(N__4289),
            .lcout(\d1.trans_up_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI5QJP_11_LC_8_10_6 .C_ON=1'b0;
    defparam \d1.count_RNI5QJP_11_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI5QJP_11_LC_8_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.count_RNI5QJP_11_LC_8_10_6  (
            .in0(N__4202),
            .in1(N__3978),
            .in2(N__4591),
            .in3(N__3527),
            .lcout(\d1.trans_up_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_RNIKI1C_LC_8_10_7 .C_ON=1'b0;
    defparam \d1.sync_1_RNIKI1C_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \d1.sync_1_RNIKI1C_LC_8_10_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \d1.sync_1_RNIKI1C_LC_8_10_7  (
            .in0(N__3528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3513),
            .lcout(\d1.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_1_LC_8_11_1 .C_ON=1'b0;
    defparam \d1.count_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \d1.count_1_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \d1.count_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__3984),
            .in2(_gnd_net_),
            .in3(N__4008),
            .lcout(\d1.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4794),
            .ce(),
            .sr(N__4506));
    defparam \d1.count_0_LC_8_11_5 .C_ON=1'b0;
    defparam \d1.count_0_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \d1.count_0_LC_8_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \d1.count_0_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3983),
            .lcout(\d1.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4794),
            .ce(),
            .sr(N__4506));
    defparam \p.count_RNIL0L01_15_LC_8_12_1 .C_ON=1'b0;
    defparam \p.count_RNIL0L01_15_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \p.count_RNIL0L01_15_LC_8_12_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \p.count_RNIL0L01_15_LC_8_12_1  (
            .in0(N__3938),
            .in1(N__3920),
            .in2(N__3900),
            .in3(N__3875),
            .lcout(\p.count10_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.count_RNIFQK01_12_LC_8_12_2 .C_ON=1'b0;
    defparam \p.count_RNIFQK01_12_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \p.count_RNIFQK01_12_LC_8_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \p.count_RNIFQK01_12_LC_8_12_2  (
            .in0(N__3854),
            .in1(N__3833),
            .in2(N__3814),
            .in3(N__3788),
            .lcout(\p.count10_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.count_RNICNK01_10_LC_8_12_5 .C_ON=1'b0;
    defparam \p.count_RNICNK01_10_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \p.count_RNICNK01_10_LC_8_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \p.count_RNICNK01_10_LC_8_12_5  (
            .in0(N__3767),
            .in1(N__3746),
            .in2(N__3727),
            .in3(N__3701),
            .lcout(),
            .ltout(\p.count10_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.count_RNIIMK74_10_LC_8_12_6 .C_ON=1'b0;
    defparam \p.count_RNIIMK74_10_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \p.count_RNIIMK74_10_LC_8_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \p.count_RNIIMK74_10_LC_8_12_6  (
            .in0(N__3682),
            .in1(N__3676),
            .in2(N__3670),
            .in3(N__3601),
            .lcout(\p.count10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \p.count_RNI24M51_1_LC_8_12_7 .C_ON=1'b0;
    defparam \p.count_RNI24M51_1_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \p.count_RNI24M51_1_LC_8_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \p.count_RNI24M51_1_LC_8_12_7  (
            .in0(N__4459),
            .in1(N__3641),
            .in2(N__4488),
            .in3(N__3620),
            .lcout(\p.count10_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIE4R8_16_LC_8_14_0 .C_ON=1'b0;
    defparam \d2.count_RNIE4R8_16_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIE4R8_16_LC_8_14_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \d2.count_RNIE4R8_16_LC_8_14_0  (
            .in0(N__4870),
            .in1(N__4887),
            .in2(_gnd_net_),
            .in3(N__4731),
            .lcout(\d2.trans_up_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNI6TT21_3_LC_8_14_1 .C_ON=1'b0;
    defparam \d2.count_RNI6TT21_3_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNI6TT21_3_LC_8_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNI6TT21_3_LC_8_14_1  (
            .in0(N__4686),
            .in1(N__4701),
            .in2(N__4672),
            .in3(N__4716),
            .lcout(\d2.trans_up_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNITE8Q_10_LC_8_14_7 .C_ON=1'b0;
    defparam \d2.count_RNITE8Q_10_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNITE8Q_10_LC_8_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNITE8Q_10_LC_8_14_7  (
            .in0(N__4623),
            .in1(N__4638),
            .in2(N__4609),
            .in3(N__4653),
            .lcout(\d2.trans_up_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNI237_11_LC_8_16_5 .C_ON=1'b0;
    defparam \d2.count_RNI237_11_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNI237_11_LC_8_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNI237_11_LC_8_16_5  (
            .in0(N__4935),
            .in1(N__4950),
            .in2(N__4921),
            .in3(N__4902),
            .lcout(\d2.count_RNI237Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_0_LC_9_4_0 .C_ON=1'b0;
    defparam \d2.sync_0_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \d2.sync_0_LC_9_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d2.sync_0_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4159),
            .lcout(\d2.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4811),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_LC_9_7_3 .C_ON=1'b0;
    defparam \d2.sync_1_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \d2.sync_1_LC_9_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d2.sync_1_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4138),
            .lcout(\d2.syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4804),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_RNIMV5K_LC_9_7_6 .C_ON=1'b0;
    defparam \d2.sync_1_RNIMV5K_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \d2.sync_1_RNIMV5K_LC_9_7_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \d2.sync_1_RNIMV5K_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__4129),
            .in2(_gnd_net_),
            .in3(N__4100),
            .lcout(\d2.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_0_LC_9_8_1 .C_ON=1'b0;
    defparam \d2.count_0_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \d2.count_0_LC_9_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \d2.count_0_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4400),
            .lcout(\d2.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4801),
            .ce(),
            .sr(N__4855));
    defparam \d2.count_1_LC_9_8_7 .C_ON=1'b0;
    defparam \d2.count_1_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_1_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \d2.count_1_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__4374),
            .in2(_gnd_net_),
            .in3(N__4401),
            .lcout(\d2.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4801),
            .ce(),
            .sr(N__4855));
    defparam \d1.un3_count_cry_1_c_LC_9_9_0 .C_ON=1'b1;
    defparam \d1.un3_count_cry_1_c_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \d1.un3_count_cry_1_c_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d1.un3_count_cry_1_c_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__4009),
            .in2(N__3988),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\d1.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_2_LC_9_9_1 .C_ON=1'b1;
    defparam \d1.count_2_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \d1.count_2_LC_9_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_2_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__3958),
            .in2(_gnd_net_),
            .in3(N__3946),
            .lcout(\d1.countZ0Z_2 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_1 ),
            .carryout(\d1.un3_count_cry_2 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_3_LC_9_9_2 .C_ON=1'b1;
    defparam \d1.count_3_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \d1.count_3_LC_9_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_3_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__4354),
            .in2(_gnd_net_),
            .in3(N__4342),
            .lcout(\d1.countZ0Z_3 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_2 ),
            .carryout(\d1.un3_count_cry_3 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_4_LC_9_9_3 .C_ON=1'b1;
    defparam \d1.count_4_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \d1.count_4_LC_9_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_4_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__4339),
            .in2(_gnd_net_),
            .in3(N__4327),
            .lcout(\d1.countZ0Z_4 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_3 ),
            .carryout(\d1.un3_count_cry_4 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_5_LC_9_9_4 .C_ON=1'b1;
    defparam \d1.count_5_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \d1.count_5_LC_9_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_5_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__4324),
            .in2(_gnd_net_),
            .in3(N__4312),
            .lcout(\d1.countZ0Z_5 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_4 ),
            .carryout(\d1.un3_count_cry_5 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_6_LC_9_9_5 .C_ON=1'b1;
    defparam \d1.count_6_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \d1.count_6_LC_9_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_6_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__4308),
            .in2(_gnd_net_),
            .in3(N__4294),
            .lcout(\d1.countZ0Z_6 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_5 ),
            .carryout(\d1.un3_count_cry_6 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_7_LC_9_9_6 .C_ON=1'b1;
    defparam \d1.count_7_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \d1.count_7_LC_9_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_7_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__4291),
            .in2(_gnd_net_),
            .in3(N__4276),
            .lcout(\d1.countZ0Z_7 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_6 ),
            .carryout(\d1.un3_count_cry_7 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_8_LC_9_9_7 .C_ON=1'b1;
    defparam \d1.count_8_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \d1.count_8_LC_9_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_8_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__4273),
            .in2(_gnd_net_),
            .in3(N__4255),
            .lcout(\d1.countZ0Z_8 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_7 ),
            .carryout(\d1.un3_count_cry_8 ),
            .clk(N__4799),
            .ce(),
            .sr(N__4507));
    defparam \d1.count_9_LC_9_10_0 .C_ON=1'b1;
    defparam \d1.count_9_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \d1.count_9_LC_9_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_9_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__4252),
            .in2(_gnd_net_),
            .in3(N__4237),
            .lcout(\d1.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\d1.un3_count_cry_9 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_10_LC_9_10_1 .C_ON=1'b1;
    defparam \d1.count_10_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \d1.count_10_LC_9_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_10_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__4229),
            .in2(_gnd_net_),
            .in3(N__4207),
            .lcout(\d1.countZ0Z_10 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_9 ),
            .carryout(\d1.un3_count_cry_10 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_11_LC_9_10_2 .C_ON=1'b1;
    defparam \d1.count_11_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \d1.count_11_LC_9_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_11_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__4204),
            .in2(_gnd_net_),
            .in3(N__4189),
            .lcout(\d1.countZ0Z_11 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_10 ),
            .carryout(\d1.un3_count_cry_11 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_12_LC_9_10_3 .C_ON=1'b1;
    defparam \d1.count_12_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \d1.count_12_LC_9_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_12_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__4590),
            .in2(_gnd_net_),
            .in3(N__4573),
            .lcout(\d1.countZ0Z_12 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_11 ),
            .carryout(\d1.un3_count_cry_12 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_13_LC_9_10_4 .C_ON=1'b1;
    defparam \d1.count_13_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \d1.count_13_LC_9_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_13_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__4570),
            .in2(_gnd_net_),
            .in3(N__4558),
            .lcout(\d1.countZ0Z_13 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_12 ),
            .carryout(\d1.un3_count_cry_13 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_14_LC_9_10_5 .C_ON=1'b1;
    defparam \d1.count_14_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \d1.count_14_LC_9_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_14_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__4555),
            .in2(_gnd_net_),
            .in3(N__4543),
            .lcout(\d1.countZ0Z_14 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_13 ),
            .carryout(\d1.un3_count_cry_14 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_15_LC_9_10_6 .C_ON=1'b1;
    defparam \d1.count_15_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \d1.count_15_LC_9_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_15_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__4540),
            .in2(_gnd_net_),
            .in3(N__4528),
            .lcout(\d1.countZ0Z_15 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_14 ),
            .carryout(\d1.un3_count_cry_15 ),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \d1.count_16_LC_9_10_7 .C_ON=1'b0;
    defparam \d1.count_16_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \d1.count_16_LC_9_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d1.count_16_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__4521),
            .in2(_gnd_net_),
            .in3(N__4525),
            .lcout(\d1.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4795),
            .ce(),
            .sr(N__4505));
    defparam \p.count_1_LC_9_12_3 .C_ON=1'b0;
    defparam \p.count_1_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \p.count_1_LC_9_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \p.count_1_LC_9_12_3  (
            .in0(N__4464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4487),
            .lcout(\p.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4791),
            .ce(N__4430),
            .sr(_gnd_net_));
    defparam \p.count_0_LC_9_12_4 .C_ON=1'b0;
    defparam \p.count_0_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \p.count_0_LC_9_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \p.count_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4463),
            .lcout(\p.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4791),
            .ce(N__4430),
            .sr(_gnd_net_));
    defparam \d2.un3_count_cry_1_c_LC_9_14_0 .C_ON=1'b1;
    defparam \d2.un3_count_cry_1_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \d2.un3_count_cry_1_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d2.un3_count_cry_1_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__4402),
            .in2(N__4378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\d2.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_2_LC_9_14_1 .C_ON=1'b1;
    defparam \d2.count_2_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \d2.count_2_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_2_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__4732),
            .in2(_gnd_net_),
            .in3(N__4720),
            .lcout(\d2.countZ0Z_2 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_1 ),
            .carryout(\d2.un3_count_cry_2 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_3_LC_9_14_2 .C_ON=1'b1;
    defparam \d2.count_3_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \d2.count_3_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_3_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__4717),
            .in2(_gnd_net_),
            .in3(N__4705),
            .lcout(\d2.countZ0Z_3 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_2 ),
            .carryout(\d2.un3_count_cry_3 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_4_LC_9_14_3 .C_ON=1'b1;
    defparam \d2.count_4_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \d2.count_4_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_4_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__4702),
            .in2(_gnd_net_),
            .in3(N__4690),
            .lcout(\d2.countZ0Z_4 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_3 ),
            .carryout(\d2.un3_count_cry_4 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_5_LC_9_14_4 .C_ON=1'b1;
    defparam \d2.count_5_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \d2.count_5_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_5_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__4687),
            .in2(_gnd_net_),
            .in3(N__4675),
            .lcout(\d2.countZ0Z_5 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_4 ),
            .carryout(\d2.un3_count_cry_5 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_6_LC_9_14_5 .C_ON=1'b1;
    defparam \d2.count_6_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \d2.count_6_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_6_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__4671),
            .in2(_gnd_net_),
            .in3(N__4657),
            .lcout(\d2.countZ0Z_6 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_5 ),
            .carryout(\d2.un3_count_cry_6 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_7_LC_9_14_6 .C_ON=1'b1;
    defparam \d2.count_7_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \d2.count_7_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_7_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__4654),
            .in2(_gnd_net_),
            .in3(N__4642),
            .lcout(\d2.countZ0Z_7 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_6 ),
            .carryout(\d2.un3_count_cry_7 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_8_LC_9_14_7 .C_ON=1'b1;
    defparam \d2.count_8_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_8_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_8_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__4639),
            .in2(_gnd_net_),
            .in3(N__4627),
            .lcout(\d2.countZ0Z_8 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_7 ),
            .carryout(\d2.un3_count_cry_8 ),
            .clk(N__4790),
            .ce(),
            .sr(N__4854));
    defparam \d2.count_9_LC_9_15_0 .C_ON=1'b1;
    defparam \d2.count_9_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \d2.count_9_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_9_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__4624),
            .in2(_gnd_net_),
            .in3(N__4612),
            .lcout(\d2.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\d2.un3_count_cry_9 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_10_LC_9_15_1 .C_ON=1'b1;
    defparam \d2.count_10_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \d2.count_10_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_10_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__4605),
            .in2(_gnd_net_),
            .in3(N__4954),
            .lcout(\d2.countZ0Z_10 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_9 ),
            .carryout(\d2.un3_count_cry_10 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_11_LC_9_15_2 .C_ON=1'b1;
    defparam \d2.count_11_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \d2.count_11_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_11_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__4951),
            .in2(_gnd_net_),
            .in3(N__4939),
            .lcout(\d2.countZ0Z_11 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_10 ),
            .carryout(\d2.un3_count_cry_11 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_12_LC_9_15_3 .C_ON=1'b1;
    defparam \d2.count_12_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \d2.count_12_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_12_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__4936),
            .in2(_gnd_net_),
            .in3(N__4924),
            .lcout(\d2.countZ0Z_12 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_11 ),
            .carryout(\d2.un3_count_cry_12 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_13_LC_9_15_4 .C_ON=1'b1;
    defparam \d2.count_13_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \d2.count_13_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_13_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__4920),
            .in2(_gnd_net_),
            .in3(N__4906),
            .lcout(\d2.countZ0Z_13 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_12 ),
            .carryout(\d2.un3_count_cry_13 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_14_LC_9_15_5 .C_ON=1'b1;
    defparam \d2.count_14_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \d2.count_14_LC_9_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_14_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__4903),
            .in2(_gnd_net_),
            .in3(N__4891),
            .lcout(\d2.countZ0Z_14 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_13 ),
            .carryout(\d2.un3_count_cry_14 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_15_LC_9_15_6 .C_ON=1'b1;
    defparam \d2.count_15_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \d2.count_15_LC_9_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_15_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__4888),
            .in2(_gnd_net_),
            .in3(N__4876),
            .lcout(\d2.countZ0Z_15 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_14 ),
            .carryout(\d2.un3_count_cry_15 ),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d2.count_16_LC_9_15_7 .C_ON=1'b0;
    defparam \d2.count_16_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_16_LC_9_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d2.count_16_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__4869),
            .in2(_gnd_net_),
            .in3(N__4873),
            .lcout(\d2.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4789),
            .ce(),
            .sr(N__4853));
    defparam \d1.sync_0_LC_10_9_3 .C_ON=1'b0;
    defparam \d1.sync_0_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \d1.sync_0_LC_10_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d1.sync_0_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4840),
            .lcout(\d1.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(_gnd_net_));
endmodule // servo_tester
