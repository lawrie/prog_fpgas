-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Dec 23 2017 18:12:09

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "servo_tester" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of servo_tester
entity servo_tester is
port (
    switch_up : in std_logic;
    switch_dn : in std_logic;
    CONTROL_PIN : out std_logic;
    CLK : in std_logic);
end servo_tester;

-- Architecture of servo_tester
-- View name is \INTERFACE\
architecture \INTERFACE\ of servo_tester is

signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \p.prescaler12_0\ : std_logic;
signal \p.prescaler12_1\ : std_logic;
signal \p.prescaler12_2\ : std_logic;
signal \p.prescaler12_3\ : std_logic;
signal \p.prescaler12_4\ : std_logic;
signal \p.prescaler12_5\ : std_logic;
signal \p.prescaler12\ : std_logic;
signal \p.prescaler12_THRU_CO\ : std_logic;
signal \p.prescaler12_4_and\ : std_logic;
signal \p.prescaler12_2_and\ : std_logic;
signal \p.prescaler12_6_and\ : std_logic;
signal \p.prescaler12_5_and\ : std_logic;
signal \p.prescaler12_3_and\ : std_logic;
signal \p.prescaler12_1_and\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \p.prescalerZ0Z_2\ : std_logic;
signal \p.prescaler_1_cry_1_THRU_CO\ : std_logic;
signal \p.prescaler_1_cry_1\ : std_logic;
signal \p.prescalerZ0Z_3\ : std_logic;
signal \p.prescaler_1_cry_2\ : std_logic;
signal \p.prescalerZ0Z_4\ : std_logic;
signal \p.prescaler_1_cry_3\ : std_logic;
signal \p.prescaler_1_cry_4\ : std_logic;
signal \p.prescaler_1_cry_5\ : std_logic;
signal \p.prescalerZ0Z_7\ : std_logic;
signal \p.prescaler_1_cry_6\ : std_logic;
signal \p.prescalerZ0Z_8\ : std_logic;
signal \p.prescaler_1_cry_7\ : std_logic;
signal \p.prescaler_1_cry_8\ : std_logic;
signal \p.prescalerZ0Z_9\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \p.prescalerZ0Z_10\ : std_logic;
signal \p.prescaler_1_cry_9\ : std_logic;
signal \p.prescalerZ0Z_11\ : std_logic;
signal \p.prescaler_1_cry_10\ : std_logic;
signal \p.prescalerZ0Z_12\ : std_logic;
signal \p.prescaler_1_cry_11\ : std_logic;
signal \p.prescalerZ0Z_13\ : std_logic;
signal \p.prescaler_1_cry_12\ : std_logic;
signal \p.prescalerZ0Z_14\ : std_logic;
signal \p.prescaler_1_cry_13\ : std_logic;
signal \p.prescalerZ0Z_15\ : std_logic;
signal \p.prescaler_1_cry_14\ : std_logic;
signal \p.prescalerZ0Z_16\ : std_logic;
signal \p.prescaler_1_cry_15\ : std_logic;
signal \p.prescaler_1_cry_16\ : std_logic;
signal \p.prescalerZ0Z_17\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \p.prescalerZ0Z_18\ : std_logic;
signal \p.prescaler_1_cry_17\ : std_logic;
signal \p.prescalerZ0Z_19\ : std_logic;
signal \p.prescaler_1_cry_18\ : std_logic;
signal \p.prescalerZ0Z_20\ : std_logic;
signal \p.prescaler_1_cry_19\ : std_logic;
signal \p.prescalerZ0Z_21\ : std_logic;
signal \p.prescaler_1_cry_20\ : std_logic;
signal \p.prescalerZ0Z_22\ : std_logic;
signal \p.prescaler_1_cry_21\ : std_logic;
signal \p.prescalerZ0Z_23\ : std_logic;
signal \p.prescaler_1_cry_22\ : std_logic;
signal \p.prescalerZ0Z_24\ : std_logic;
signal \p.prescaler_1_cry_23\ : std_logic;
signal \p.prescaler_1_cry_24\ : std_logic;
signal \p.prescalerZ0Z_25\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \p.prescaler_1_cry_25\ : std_logic;
signal \p.prescalerZ0Z_26\ : std_logic;
signal \p.prescaler12_0_and\ : std_logic;
signal \p.prescaler_1_cry_5_THRU_CO\ : std_logic;
signal \p.prescalerZ0Z_6\ : std_logic;
signal \p.prescaler_1_cry_4_THRU_CO\ : std_logic;
signal \p.prescalerZ0Z_5\ : std_logic;
signal \p.prescalerZ0Z_0\ : std_logic;
signal \p.prescalerZ0Z_1\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \state_RNIPC4P3\ : std_logic;
signal un1_pulse_len_cry_2 : std_logic;
signal un1_pulse_len_cry_3 : std_logic;
signal un1_pulse_len_cry_4 : std_logic;
signal un1_pulse_len_cry_5 : std_logic;
signal un1_pulse_len_cry_6 : std_logic;
signal \state_RNIPC4P3_6\ : std_logic;
signal un1_pulse_len_cry_7 : std_logic;
signal un1_pulse_len_cry_8 : std_logic;
signal un1_pulse_len_cry_9 : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal un1_pulse_len_cry_10 : std_logic;
signal un1_pulse_len_cry_11 : std_logic;
signal un1_pulse_len_cry_12 : std_logic;
signal un1_pulse_len_cry_13 : std_logic;
signal un1_pulse_len_cry_14 : std_logic;
signal \state_RNIPC4P3_4\ : std_logic;
signal \state_RNIPC4P3_7\ : std_logic;
signal \p.count_i_2\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \pulse_lenZ0Z_3\ : std_logic;
signal \p.count_i_3\ : std_logic;
signal \p.CONTROL_PIN_2_cry_2\ : std_logic;
signal \pulse_lenZ0Z_4\ : std_logic;
signal \p.count_i_4\ : std_logic;
signal \p.CONTROL_PIN_2_cry_3\ : std_logic;
signal \pulse_lenZ0Z_5\ : std_logic;
signal \p.count_i_5\ : std_logic;
signal \p.CONTROL_PIN_2_cry_4\ : std_logic;
signal \pulse_lenZ0Z_6\ : std_logic;
signal \p.count_i_6\ : std_logic;
signal \p.CONTROL_PIN_2_cry_5\ : std_logic;
signal \pulse_lenZ0Z_7\ : std_logic;
signal \p.count_i_7\ : std_logic;
signal \p.CONTROL_PIN_2_cry_6\ : std_logic;
signal \pulse_lenZ0Z_8\ : std_logic;
signal \p.count_i_8\ : std_logic;
signal \p.CONTROL_PIN_2_cry_7\ : std_logic;
signal \pulse_lenZ0Z_9\ : std_logic;
signal \p.count_i_9\ : std_logic;
signal \p.CONTROL_PIN_2_cry_8\ : std_logic;
signal \p.CONTROL_PIN_2_cry_9\ : std_logic;
signal \pulse_lenZ0Z_10\ : std_logic;
signal \p.count_i_10\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \pulse_lenZ0Z_11\ : std_logic;
signal \p.count_i_11\ : std_logic;
signal \p.CONTROL_PIN_2_cry_10\ : std_logic;
signal \pulse_lenZ0Z_12\ : std_logic;
signal \p.count_i_12\ : std_logic;
signal \p.CONTROL_PIN_2_cry_11\ : std_logic;
signal \pulse_lenZ0Z_13\ : std_logic;
signal \p.count_i_13\ : std_logic;
signal \p.CONTROL_PIN_2_cry_12\ : std_logic;
signal \pulse_lenZ0Z_14\ : std_logic;
signal \p.count_i_14\ : std_logic;
signal \p.CONTROL_PIN_2_cry_13\ : std_logic;
signal \pulse_lenZ0Z_15\ : std_logic;
signal \p.count_i_15\ : std_logic;
signal \p.CONTROL_PIN_2_cry_14\ : std_logic;
signal \p.CONTROL_PIN_2\ : std_logic;
signal \CONTROL_PIN_c\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \p.count_1_cry_1\ : std_logic;
signal \p.count_1_cry_2\ : std_logic;
signal \p.count_1_cry_3\ : std_logic;
signal \p.count_1_cry_4\ : std_logic;
signal \p.count_1_cry_5\ : std_logic;
signal \p.count_1_cry_6\ : std_logic;
signal \p.count_1_cry_7\ : std_logic;
signal \p.count_1_cry_8\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \p.count_1_cry_9\ : std_logic;
signal \p.count_1_cry_10\ : std_logic;
signal \p.count_1_cry_11\ : std_logic;
signal \p.count_1_cry_12\ : std_logic;
signal \p.count_1_cry_13\ : std_logic;
signal \p.count_1_cry_14\ : std_logic;
signal \state_RNIPC4P3_0\ : std_logic;
signal \state_RNIPC4P3_2\ : std_logic;
signal \d2.trans_up_1_12_cascade_\ : std_logic;
signal \d2.trans_up_1_sx_cascade_\ : std_logic;
signal \d2_trans_up_1_cascade_\ : std_logic;
signal \pulse_lenZ0Z_2\ : std_logic;
signal \s_dn_i_cascade_\ : std_logic;
signal \un1_pulse_len_cry_2_c_RNOZ0\ : std_logic;
signal \state_RNIPC4P3_3\ : std_logic;
signal \state_RNIU5D07\ : std_logic;
signal \state_RNIPC4P3_1\ : std_logic;
signal \state_RNIPC4P3_8\ : std_logic;
signal d2_trans_up_1 : std_logic;
signal \state_RNIPC4P3_5\ : std_logic;
signal \d1.count_RNI2PCEZ0Z_3_cascade_\ : std_logic;
signal \d1.trans_up_1_14_cascade_\ : std_logic;
signal s_up : std_logic;
signal \s_up_cascade_\ : std_logic;
signal s_dn_i : std_logic;
signal \state_RNIU5D07_0\ : std_logic;
signal \d1.trans_up_1_11\ : std_logic;
signal \d1.trans_up_1_13_sx_cascade_\ : std_logic;
signal \d1.trans_up_1_14\ : std_logic;
signal \d1.trans_up_1_13_cascade_\ : std_logic;
signal \d1.trans_up_1_12\ : std_logic;
signal \d1.trans_up_1_9\ : std_logic;
signal \d1.trans_up_sx\ : std_logic;
signal \d1.stateZ0\ : std_logic;
signal \d1.syncZ0Z_1\ : std_logic;
signal \d1.idle_i\ : std_logic;
signal \p.countZ0Z_14\ : std_logic;
signal \p.countZ0Z_8\ : std_logic;
signal \p.countZ0Z_15\ : std_logic;
signal \p.countZ0Z_6\ : std_logic;
signal \p.countZ0Z_12\ : std_logic;
signal \p.countZ0Z_7\ : std_logic;
signal \p.countZ0Z_13\ : std_logic;
signal \p.countZ0Z_5\ : std_logic;
signal \p.countZ0Z_10\ : std_logic;
signal \p.countZ0Z_9\ : std_logic;
signal \p.countZ0Z_11\ : std_logic;
signal \p.countZ0Z_4\ : std_logic;
signal \p.count10_11\ : std_logic;
signal \p.count10_10\ : std_logic;
signal \p.count10_8_cascade_\ : std_logic;
signal \p.count10\ : std_logic;
signal \p.countZ0Z_3\ : std_logic;
signal \p.countZ0Z_2\ : std_logic;
signal \p.count10_9\ : std_logic;
signal \d2.trans_up_1_11\ : std_logic;
signal \d2.trans_up_1_10\ : std_logic;
signal \d2.trans_up_1_9\ : std_logic;
signal \d2.count_RNI237Z0Z_11\ : std_logic;
signal switch_dn_c : std_logic;
signal \d2.syncZ0Z_0\ : std_logic;
signal \d2.syncZ0Z_1\ : std_logic;
signal d2_state : std_logic;
signal \d2.idle_i\ : std_logic;
signal \d1.countZ0Z_1\ : std_logic;
signal \d1.countZ0Z_0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \d1.countZ0Z_2\ : std_logic;
signal \d1.un3_count_cry_1\ : std_logic;
signal \d1.countZ0Z_3\ : std_logic;
signal \d1.un3_count_cry_2\ : std_logic;
signal \d1.countZ0Z_4\ : std_logic;
signal \d1.un3_count_cry_3\ : std_logic;
signal \d1.countZ0Z_5\ : std_logic;
signal \d1.un3_count_cry_4\ : std_logic;
signal \d1.countZ0Z_6\ : std_logic;
signal \d1.un3_count_cry_5\ : std_logic;
signal \d1.countZ0Z_7\ : std_logic;
signal \d1.un3_count_cry_6\ : std_logic;
signal \d1.countZ0Z_8\ : std_logic;
signal \d1.un3_count_cry_7\ : std_logic;
signal \d1.un3_count_cry_8\ : std_logic;
signal \d1.countZ0Z_9\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \d1.countZ0Z_10\ : std_logic;
signal \d1.un3_count_cry_9\ : std_logic;
signal \d1.countZ0Z_11\ : std_logic;
signal \d1.un3_count_cry_10\ : std_logic;
signal \d1.countZ0Z_12\ : std_logic;
signal \d1.un3_count_cry_11\ : std_logic;
signal \d1.countZ0Z_13\ : std_logic;
signal \d1.un3_count_cry_12\ : std_logic;
signal \d1.countZ0Z_14\ : std_logic;
signal \d1.un3_count_cry_13\ : std_logic;
signal \d1.countZ0Z_15\ : std_logic;
signal \d1.un3_count_cry_14\ : std_logic;
signal \d1.un3_count_cry_15\ : std_logic;
signal \d1.countZ0Z_16\ : std_logic;
signal \d1.idle_i_g\ : std_logic;
signal \p.countZ0Z_1\ : std_logic;
signal \p.countZ0Z_0\ : std_logic;
signal \p.prescaler12_g\ : std_logic;
signal \d2.countZ0Z_0\ : std_logic;
signal \d2.countZ0Z_1\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \d2.countZ0Z_2\ : std_logic;
signal \d2.un3_count_cry_1\ : std_logic;
signal \d2.countZ0Z_3\ : std_logic;
signal \d2.un3_count_cry_2\ : std_logic;
signal \d2.countZ0Z_4\ : std_logic;
signal \d2.un3_count_cry_3\ : std_logic;
signal \d2.countZ0Z_5\ : std_logic;
signal \d2.un3_count_cry_4\ : std_logic;
signal \d2.countZ0Z_6\ : std_logic;
signal \d2.un3_count_cry_5\ : std_logic;
signal \d2.countZ0Z_7\ : std_logic;
signal \d2.un3_count_cry_6\ : std_logic;
signal \d2.countZ0Z_8\ : std_logic;
signal \d2.un3_count_cry_7\ : std_logic;
signal \d2.un3_count_cry_8\ : std_logic;
signal \d2.countZ0Z_9\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \d2.countZ0Z_10\ : std_logic;
signal \d2.un3_count_cry_9\ : std_logic;
signal \d2.countZ0Z_11\ : std_logic;
signal \d2.un3_count_cry_10\ : std_logic;
signal \d2.countZ0Z_12\ : std_logic;
signal \d2.un3_count_cry_11\ : std_logic;
signal \d2.countZ0Z_13\ : std_logic;
signal \d2.un3_count_cry_12\ : std_logic;
signal \d2.countZ0Z_14\ : std_logic;
signal \d2.un3_count_cry_13\ : std_logic;
signal \d2.countZ0Z_15\ : std_logic;
signal \d2.un3_count_cry_14\ : std_logic;
signal \d2.un3_count_cry_15\ : std_logic;
signal \d2.countZ0Z_16\ : std_logic;
signal \d2.idle_i_g\ : std_logic;
signal switch_up_c : std_logic;
signal \d1.syncZ0Z_0\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \CONTROL_PIN_wire\ : std_logic;
signal switch_dn_wire : std_logic;
signal switch_up_wire : std_logic;

begin
    \CLK_wire\ <= CLK;
    CONTROL_PIN <= \CONTROL_PIN_wire\;
    switch_dn_wire <= switch_dn;
    switch_up_wire <= switch_up;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5000\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5002\,
            DIN => \N__5001\,
            DOUT => \N__5000\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5002\,
            PADOUT => \N__5001\,
            PADIN => \N__5000\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CONTROL_PIN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4991\,
            DIN => \N__4990\,
            DOUT => \N__4989\,
            PACKAGEPIN => \CONTROL_PIN_wire\
        );

    \CONTROL_PIN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4991\,
            PADOUT => \N__4990\,
            PADIN => \N__4989\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3235\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_dn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4982\,
            DIN => \N__4981\,
            DOUT => \N__4980\,
            PACKAGEPIN => switch_dn_wire
        );

    \switch_dn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4982\,
            PADOUT => \N__4981\,
            PADIN => \N__4980\,
            CLOCKENABLE => 'H',
            DIN0 => switch_dn_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \switch_up_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4973\,
            DIN => \N__4972\,
            DOUT => \N__4971\,
            PACKAGEPIN => switch_up_wire
        );

    \switch_up_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4973\,
            PADOUT => \N__4972\,
            PADIN => \N__4971\,
            CLOCKENABLE => 'H',
            DIN0 => switch_up_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1092\ : InMux
    port map (
            O => \N__4954\,
            I => \d2.un3_count_cry_9\
        );

    \I__1091\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4947\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4944\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4947\,
            I => \d2.countZ0Z_11\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4944\,
            I => \d2.countZ0Z_11\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4939\,
            I => \d2.un3_count_cry_10\
        );

    \I__1086\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4932\
        );

    \I__1085\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4929\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__4932\,
            I => \d2.countZ0Z_12\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__4929\,
            I => \d2.countZ0Z_12\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4924\,
            I => \d2.un3_count_cry_11\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__4921\,
            I => \N__4917\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4914\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4911\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4914\,
            I => \d2.countZ0Z_13\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4911\,
            I => \d2.countZ0Z_13\
        );

    \I__1076\ : InMux
    port map (
            O => \N__4906\,
            I => \d2.un3_count_cry_12\
        );

    \I__1075\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4899\
        );

    \I__1074\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4896\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__4899\,
            I => \d2.countZ0Z_14\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4896\,
            I => \d2.countZ0Z_14\
        );

    \I__1071\ : InMux
    port map (
            O => \N__4891\,
            I => \d2.un3_count_cry_13\
        );

    \I__1070\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4884\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4881\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4884\,
            I => \d2.countZ0Z_15\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__4881\,
            I => \d2.countZ0Z_15\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4876\,
            I => \d2.un3_count_cry_14\
        );

    \I__1065\ : InMux
    port map (
            O => \N__4873\,
            I => \d2.un3_count_cry_15\
        );

    \I__1064\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4866\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4863\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__4866\,
            I => \N__4860\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4863\,
            I => \d2.countZ0Z_16\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__4860\,
            I => \d2.countZ0Z_16\
        );

    \I__1059\ : SRMux
    port map (
            O => \N__4855\,
            I => \N__4846\
        );

    \I__1058\ : SRMux
    port map (
            O => \N__4854\,
            I => \N__4846\
        );

    \I__1057\ : SRMux
    port map (
            O => \N__4853\,
            I => \N__4846\
        );

    \I__1056\ : GlobalMux
    port map (
            O => \N__4846\,
            I => \N__4843\
        );

    \I__1055\ : gio2CtrlBuf
    port map (
            O => \N__4843\,
            I => \d2.idle_i_g\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__1052\ : Span12Mux_h
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__1051\ : Span12Mux_v
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__1050\ : Span12Mux_h
    port map (
            O => \N__4828\,
            I => \N__4825\
        );

    \I__1049\ : Odrv12
    port map (
            O => \N__4825\,
            I => switch_up_c
        );

    \I__1048\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__4816\,
            I => \d1.syncZ0Z_0\
        );

    \I__1045\ : ClkMux
    port map (
            O => \N__4813\,
            I => \N__4738\
        );

    \I__1044\ : ClkMux
    port map (
            O => \N__4812\,
            I => \N__4738\
        );

    \I__1043\ : ClkMux
    port map (
            O => \N__4811\,
            I => \N__4738\
        );

    \I__1042\ : ClkMux
    port map (
            O => \N__4810\,
            I => \N__4738\
        );

    \I__1041\ : ClkMux
    port map (
            O => \N__4809\,
            I => \N__4738\
        );

    \I__1040\ : ClkMux
    port map (
            O => \N__4808\,
            I => \N__4738\
        );

    \I__1039\ : ClkMux
    port map (
            O => \N__4807\,
            I => \N__4738\
        );

    \I__1038\ : ClkMux
    port map (
            O => \N__4806\,
            I => \N__4738\
        );

    \I__1037\ : ClkMux
    port map (
            O => \N__4805\,
            I => \N__4738\
        );

    \I__1036\ : ClkMux
    port map (
            O => \N__4804\,
            I => \N__4738\
        );

    \I__1035\ : ClkMux
    port map (
            O => \N__4803\,
            I => \N__4738\
        );

    \I__1034\ : ClkMux
    port map (
            O => \N__4802\,
            I => \N__4738\
        );

    \I__1033\ : ClkMux
    port map (
            O => \N__4801\,
            I => \N__4738\
        );

    \I__1032\ : ClkMux
    port map (
            O => \N__4800\,
            I => \N__4738\
        );

    \I__1031\ : ClkMux
    port map (
            O => \N__4799\,
            I => \N__4738\
        );

    \I__1030\ : ClkMux
    port map (
            O => \N__4798\,
            I => \N__4738\
        );

    \I__1029\ : ClkMux
    port map (
            O => \N__4797\,
            I => \N__4738\
        );

    \I__1028\ : ClkMux
    port map (
            O => \N__4796\,
            I => \N__4738\
        );

    \I__1027\ : ClkMux
    port map (
            O => \N__4795\,
            I => \N__4738\
        );

    \I__1026\ : ClkMux
    port map (
            O => \N__4794\,
            I => \N__4738\
        );

    \I__1025\ : ClkMux
    port map (
            O => \N__4793\,
            I => \N__4738\
        );

    \I__1024\ : ClkMux
    port map (
            O => \N__4792\,
            I => \N__4738\
        );

    \I__1023\ : ClkMux
    port map (
            O => \N__4791\,
            I => \N__4738\
        );

    \I__1022\ : ClkMux
    port map (
            O => \N__4790\,
            I => \N__4738\
        );

    \I__1021\ : ClkMux
    port map (
            O => \N__4789\,
            I => \N__4738\
        );

    \I__1020\ : GlobalMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__1019\ : gio2CtrlBuf
    port map (
            O => \N__4735\,
            I => \CLK_c_g\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4728\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4728\,
            I => \d2.countZ0Z_2\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4725\,
            I => \d2.countZ0Z_2\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4720\,
            I => \d2.un3_count_cry_1\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4713\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4713\,
            I => \d2.countZ0Z_3\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4710\,
            I => \d2.countZ0Z_3\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4705\,
            I => \d2.un3_count_cry_2\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4698\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4695\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4698\,
            I => \d2.countZ0Z_4\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4695\,
            I => \d2.countZ0Z_4\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4690\,
            I => \d2.un3_count_cry_3\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4683\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4680\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4683\,
            I => \d2.countZ0Z_5\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4680\,
            I => \d2.countZ0Z_5\
        );

    \I__999\ : InMux
    port map (
            O => \N__4675\,
            I => \d2.un3_count_cry_4\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__4672\,
            I => \N__4668\
        );

    \I__997\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4665\
        );

    \I__996\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4662\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4665\,
            I => \d2.countZ0Z_6\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4662\,
            I => \d2.countZ0Z_6\
        );

    \I__993\ : InMux
    port map (
            O => \N__4657\,
            I => \d2.un3_count_cry_5\
        );

    \I__992\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4650\
        );

    \I__991\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4647\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4650\,
            I => \d2.countZ0Z_7\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4647\,
            I => \d2.countZ0Z_7\
        );

    \I__988\ : InMux
    port map (
            O => \N__4642\,
            I => \d2.un3_count_cry_6\
        );

    \I__987\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4635\
        );

    \I__986\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4632\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4635\,
            I => \d2.countZ0Z_8\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4632\,
            I => \d2.countZ0Z_8\
        );

    \I__983\ : InMux
    port map (
            O => \N__4627\,
            I => \d2.un3_count_cry_7\
        );

    \I__982\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4620\
        );

    \I__981\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4617\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4620\,
            I => \d2.countZ0Z_9\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4617\,
            I => \d2.countZ0Z_9\
        );

    \I__978\ : InMux
    port map (
            O => \N__4612\,
            I => \bfn_9_15_0_\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__976\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4602\
        );

    \I__975\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4599\,
            I => \d2.countZ0Z_10\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__4596\,
            I => \d2.countZ0Z_10\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__4591\,
            I => \N__4586\
        );

    \I__970\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4583\
        );

    \I__969\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4578\
        );

    \I__968\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4578\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4583\,
            I => \d1.countZ0Z_12\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4578\,
            I => \d1.countZ0Z_12\
        );

    \I__965\ : InMux
    port map (
            O => \N__4573\,
            I => \d1.un3_count_cry_11\
        );

    \I__964\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4566\
        );

    \I__963\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4566\,
            I => \d1.countZ0Z_13\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4563\,
            I => \d1.countZ0Z_13\
        );

    \I__960\ : InMux
    port map (
            O => \N__4558\,
            I => \d1.un3_count_cry_12\
        );

    \I__959\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4551\
        );

    \I__958\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4548\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4551\,
            I => \d1.countZ0Z_14\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4548\,
            I => \d1.countZ0Z_14\
        );

    \I__955\ : InMux
    port map (
            O => \N__4543\,
            I => \d1.un3_count_cry_13\
        );

    \I__954\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4536\
        );

    \I__953\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4533\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4536\,
            I => \d1.countZ0Z_15\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4533\,
            I => \d1.countZ0Z_15\
        );

    \I__950\ : InMux
    port map (
            O => \N__4528\,
            I => \d1.un3_count_cry_14\
        );

    \I__949\ : InMux
    port map (
            O => \N__4525\,
            I => \d1.un3_count_cry_15\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__4522\,
            I => \N__4518\
        );

    \I__947\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4515\
        );

    \I__946\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4512\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4515\,
            I => \d1.countZ0Z_16\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4512\,
            I => \d1.countZ0Z_16\
        );

    \I__943\ : SRMux
    port map (
            O => \N__4507\,
            I => \N__4498\
        );

    \I__942\ : SRMux
    port map (
            O => \N__4506\,
            I => \N__4498\
        );

    \I__941\ : SRMux
    port map (
            O => \N__4505\,
            I => \N__4498\
        );

    \I__940\ : GlobalMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__939\ : gio2CtrlBuf
    port map (
            O => \N__4495\,
            I => \d1.idle_i_g\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__937\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4484\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \N__4481\
        );

    \I__935\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4478\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4484\,
            I => \N__4475\
        );

    \I__933\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4472\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4478\,
            I => \p.countZ0Z_1\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__4475\,
            I => \p.countZ0Z_1\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4472\,
            I => \p.countZ0Z_1\
        );

    \I__929\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4460\
        );

    \I__928\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4454\
        );

    \I__927\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4454\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4451\
        );

    \I__925\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4448\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4454\,
            I => \p.countZ0Z_0\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__4451\,
            I => \p.countZ0Z_0\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4448\,
            I => \p.countZ0Z_0\
        );

    \I__921\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4434\
        );

    \I__920\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4434\
        );

    \I__919\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4431\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4424\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4431\,
            I => \N__4421\
        );

    \I__916\ : CEMux
    port map (
            O => \N__4430\,
            I => \N__4408\
        );

    \I__915\ : CEMux
    port map (
            O => \N__4429\,
            I => \N__4408\
        );

    \I__914\ : CEMux
    port map (
            O => \N__4428\,
            I => \N__4408\
        );

    \I__913\ : CEMux
    port map (
            O => \N__4427\,
            I => \N__4408\
        );

    \I__912\ : Glb2LocalMux
    port map (
            O => \N__4424\,
            I => \N__4408\
        );

    \I__911\ : Glb2LocalMux
    port map (
            O => \N__4421\,
            I => \N__4408\
        );

    \I__910\ : GlobalMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__909\ : gio2CtrlBuf
    port map (
            O => \N__4405\,
            I => \p.prescaler12_g\
        );

    \I__908\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4397\
        );

    \I__907\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4391\
        );

    \I__906\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4391\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4388\
        );

    \I__904\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4385\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4391\,
            I => \d2.countZ0Z_0\
        );

    \I__902\ : Odrv12
    port map (
            O => \N__4388\,
            I => \d2.countZ0Z_0\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4385\,
            I => \d2.countZ0Z_0\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4378\,
            I => \N__4375\
        );

    \I__899\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4371\
        );

    \I__898\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4367\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4371\,
            I => \N__4364\
        );

    \I__896\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4361\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4367\,
            I => \d2.countZ0Z_1\
        );

    \I__894\ : Odrv12
    port map (
            O => \N__4364\,
            I => \d2.countZ0Z_1\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4361\,
            I => \d2.countZ0Z_1\
        );

    \I__892\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4350\
        );

    \I__891\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4347\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4350\,
            I => \d1.countZ0Z_3\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4347\,
            I => \d1.countZ0Z_3\
        );

    \I__888\ : InMux
    port map (
            O => \N__4342\,
            I => \d1.un3_count_cry_2\
        );

    \I__887\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4335\
        );

    \I__886\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4332\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4335\,
            I => \d1.countZ0Z_4\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4332\,
            I => \d1.countZ0Z_4\
        );

    \I__883\ : InMux
    port map (
            O => \N__4327\,
            I => \d1.un3_count_cry_3\
        );

    \I__882\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4320\
        );

    \I__881\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4317\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4320\,
            I => \d1.countZ0Z_5\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4317\,
            I => \d1.countZ0Z_5\
        );

    \I__878\ : InMux
    port map (
            O => \N__4312\,
            I => \d1.un3_count_cry_4\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4309\,
            I => \N__4305\
        );

    \I__876\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4302\
        );

    \I__875\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4299\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4302\,
            I => \d1.countZ0Z_6\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4299\,
            I => \d1.countZ0Z_6\
        );

    \I__872\ : InMux
    port map (
            O => \N__4294\,
            I => \d1.un3_count_cry_5\
        );

    \I__871\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4286\
        );

    \I__870\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4281\
        );

    \I__869\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4281\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4286\,
            I => \d1.countZ0Z_7\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4281\,
            I => \d1.countZ0Z_7\
        );

    \I__866\ : InMux
    port map (
            O => \N__4276\,
            I => \d1.un3_count_cry_6\
        );

    \I__865\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4268\
        );

    \I__864\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4265\
        );

    \I__863\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4262\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4268\,
            I => \d1.countZ0Z_8\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4265\,
            I => \d1.countZ0Z_8\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4262\,
            I => \d1.countZ0Z_8\
        );

    \I__859\ : InMux
    port map (
            O => \N__4255\,
            I => \d1.un3_count_cry_7\
        );

    \I__858\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4247\
        );

    \I__857\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4242\
        );

    \I__856\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4242\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4247\,
            I => \d1.countZ0Z_9\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4242\,
            I => \d1.countZ0Z_9\
        );

    \I__853\ : InMux
    port map (
            O => \N__4237\,
            I => \bfn_9_10_0_\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__4234\,
            I => \N__4230\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__4233\,
            I => \N__4226\
        );

    \I__850\ : InMux
    port map (
            O => \N__4230\,
            I => \N__4223\
        );

    \I__849\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4220\
        );

    \I__848\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4217\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4223\,
            I => \N__4214\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4220\,
            I => \d1.countZ0Z_10\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4217\,
            I => \d1.countZ0Z_10\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4214\,
            I => \d1.countZ0Z_10\
        );

    \I__843\ : InMux
    port map (
            O => \N__4207\,
            I => \d1.un3_count_cry_9\
        );

    \I__842\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4199\
        );

    \I__841\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4194\
        );

    \I__840\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4194\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4199\,
            I => \d1.countZ0Z_11\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4194\,
            I => \d1.countZ0Z_11\
        );

    \I__837\ : InMux
    port map (
            O => \N__4189\,
            I => \d1.un3_count_cry_10\
        );

    \I__836\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__4177\,
            I => \d2.trans_up_1_9\
        );

    \I__832\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__830\ : Span4Mux_v
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__4162\,
            I => \d2.count_RNI237Z0Z_11\
        );

    \I__827\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__823\ : Sp12to4
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__822\ : Span12Mux_h
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__821\ : Odrv12
    port map (
            O => \N__4141\,
            I => switch_dn_c
        );

    \I__820\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__818\ : Odrv12
    port map (
            O => \N__4132\,
            I => \d2.syncZ0Z_0\
        );

    \I__817\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4125\
        );

    \I__816\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4122\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4125\,
            I => \d2.syncZ0Z_1\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4122\,
            I => \d2.syncZ0Z_1\
        );

    \I__813\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4112\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__4116\,
            I => \N__4109\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__4115\,
            I => \N__4105\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4112\,
            I => \N__4097\
        );

    \I__809\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4092\
        );

    \I__808\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4092\
        );

    \I__807\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4085\
        );

    \I__806\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4085\
        );

    \I__805\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4085\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4102\,
            I => \N__4081\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__4101\,
            I => \N__4078\
        );

    \I__802\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4070\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__4097\,
            I => \N__4063\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4092\,
            I => \N__4063\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4085\,
            I => \N__4063\
        );

    \I__798\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4060\
        );

    \I__797\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4053\
        );

    \I__796\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4053\
        );

    \I__795\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4053\
        );

    \I__794\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4050\
        );

    \I__793\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4043\
        );

    \I__792\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4043\
        );

    \I__791\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4043\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4070\,
            I => d2_state
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4063\,
            I => d2_state
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4060\,
            I => d2_state
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4053\,
            I => d2_state
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4050\,
            I => d2_state
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4043\,
            I => d2_state
        );

    \I__784\ : IoInMux
    port map (
            O => \N__4030\,
            I => \N__4027\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__782\ : Span4Mux_s1_v
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__781\ : Sp12to4
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__4018\,
            I => \N__4015\
        );

    \I__779\ : Span12Mux_v
    port map (
            O => \N__4015\,
            I => \N__4012\
        );

    \I__778\ : Odrv12
    port map (
            O => \N__4012\,
            I => \d2.idle_i\
        );

    \I__777\ : InMux
    port map (
            O => \N__4009\,
            I => \N__4005\
        );

    \I__776\ : InMux
    port map (
            O => \N__4008\,
            I => \N__4001\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__3998\
        );

    \I__774\ : InMux
    port map (
            O => \N__4004\,
            I => \N__3995\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4001\,
            I => \d1.countZ0Z_1\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__3998\,
            I => \d1.countZ0Z_1\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3995\,
            I => \d1.countZ0Z_1\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__3988\,
            I => \N__3985\
        );

    \I__769\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3980\
        );

    \I__768\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3973\
        );

    \I__767\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3973\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3970\
        );

    \I__765\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3965\
        );

    \I__764\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3965\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3973\,
            I => \d1.countZ0Z_0\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__3970\,
            I => \d1.countZ0Z_0\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3965\,
            I => \d1.countZ0Z_0\
        );

    \I__760\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3954\
        );

    \I__759\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3951\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3954\,
            I => \d1.countZ0Z_2\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3951\,
            I => \d1.countZ0Z_2\
        );

    \I__756\ : InMux
    port map (
            O => \N__3946\,
            I => \d1.un3_count_cry_1\
        );

    \I__755\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3939\
        );

    \I__754\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3935\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3939\,
            I => \N__3932\
        );

    \I__752\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3929\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3935\,
            I => \p.countZ0Z_14\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__3932\,
            I => \p.countZ0Z_14\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3929\,
            I => \p.countZ0Z_14\
        );

    \I__748\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3917\
        );

    \I__747\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3914\
        );

    \I__746\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3911\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3917\,
            I => \N__3908\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3914\,
            I => \p.countZ0Z_8\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3911\,
            I => \p.countZ0Z_8\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__3908\,
            I => \p.countZ0Z_8\
        );

    \I__741\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3896\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__3900\,
            I => \N__3893\
        );

    \I__739\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3890\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3896\,
            I => \N__3887\
        );

    \I__737\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3884\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3890\,
            I => \p.countZ0Z_15\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3887\,
            I => \p.countZ0Z_15\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3884\,
            I => \p.countZ0Z_15\
        );

    \I__733\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3872\
        );

    \I__732\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3869\
        );

    \I__731\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3866\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3863\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3869\,
            I => \p.countZ0Z_6\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3866\,
            I => \p.countZ0Z_6\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__3863\,
            I => \p.countZ0Z_6\
        );

    \I__726\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3851\
        );

    \I__725\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3848\
        );

    \I__724\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3845\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3851\,
            I => \N__3842\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3848\,
            I => \p.countZ0Z_12\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3845\,
            I => \p.countZ0Z_12\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__3842\,
            I => \p.countZ0Z_12\
        );

    \I__719\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3830\
        );

    \I__718\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3827\
        );

    \I__717\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3824\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3830\,
            I => \N__3821\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3827\,
            I => \p.countZ0Z_7\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3824\,
            I => \p.countZ0Z_7\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__3821\,
            I => \p.countZ0Z_7\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__3814\,
            I => \N__3809\
        );

    \I__711\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3806\
        );

    \I__710\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3803\
        );

    \I__709\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3800\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3806\,
            I => \N__3797\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__3803\,
            I => \p.countZ0Z_13\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3800\,
            I => \p.countZ0Z_13\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__3797\,
            I => \p.countZ0Z_13\
        );

    \I__704\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3785\
        );

    \I__703\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3782\
        );

    \I__702\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3779\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3785\,
            I => \N__3776\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3782\,
            I => \p.countZ0Z_5\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3779\,
            I => \p.countZ0Z_5\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__3776\,
            I => \p.countZ0Z_5\
        );

    \I__697\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3764\
        );

    \I__696\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3761\
        );

    \I__695\ : InMux
    port map (
            O => \N__3767\,
            I => \N__3758\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3764\,
            I => \N__3755\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3761\,
            I => \p.countZ0Z_10\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3758\,
            I => \p.countZ0Z_10\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__3755\,
            I => \p.countZ0Z_10\
        );

    \I__690\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3743\
        );

    \I__689\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3740\
        );

    \I__688\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3737\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3743\,
            I => \N__3734\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3740\,
            I => \p.countZ0Z_9\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3737\,
            I => \p.countZ0Z_9\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__3734\,
            I => \p.countZ0Z_9\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__3727\,
            I => \N__3722\
        );

    \I__682\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3719\
        );

    \I__681\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3716\
        );

    \I__680\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3713\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3710\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3716\,
            I => \p.countZ0Z_11\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3713\,
            I => \p.countZ0Z_11\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3710\,
            I => \p.countZ0Z_11\
        );

    \I__675\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3698\
        );

    \I__674\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3695\
        );

    \I__673\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3692\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3689\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3695\,
            I => \p.countZ0Z_4\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3692\,
            I => \p.countZ0Z_4\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__3689\,
            I => \p.countZ0Z_4\
        );

    \I__668\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3679\,
            I => \p.count10_11\
        );

    \I__666\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3673\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3673\,
            I => \p.count10_10\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3670\,
            I => \p.count10_8_cascade_\
        );

    \I__663\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3658\
        );

    \I__662\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3658\
        );

    \I__661\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3655\
        );

    \I__660\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3650\
        );

    \I__659\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3650\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3658\,
            I => \p.count10\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3655\,
            I => \p.count10\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3650\,
            I => \p.count10\
        );

    \I__655\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3638\
        );

    \I__654\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3635\
        );

    \I__653\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3632\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3638\,
            I => \N__3629\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3635\,
            I => \p.countZ0Z_3\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3632\,
            I => \p.countZ0Z_3\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__3629\,
            I => \p.countZ0Z_3\
        );

    \I__648\ : InMux
    port map (
            O => \N__3622\,
            I => \N__3617\
        );

    \I__647\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3614\
        );

    \I__646\ : InMux
    port map (
            O => \N__3620\,
            I => \N__3611\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3617\,
            I => \N__3608\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3614\,
            I => \p.countZ0Z_2\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3611\,
            I => \p.countZ0Z_2\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__3608\,
            I => \p.countZ0Z_2\
        );

    \I__641\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3598\,
            I => \p.count10_9\
        );

    \I__639\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__3589\,
            I => \N__3586\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__3586\,
            I => \d2.trans_up_1_11\
        );

    \I__635\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3580\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__3577\,
            I => \N__3574\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3574\,
            I => \d2.trans_up_1_10\
        );

    \I__631\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3568\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3568\,
            I => \d1.trans_up_1_11\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3565\,
            I => \d1.trans_up_1_13_sx_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3559\,
            I => \d1.trans_up_1_14\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__3556\,
            I => \d1.trans_up_1_13_cascade_\
        );

    \I__625\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3549\
        );

    \I__624\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3546\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3549\,
            I => \d1.trans_up_1_12\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3546\,
            I => \d1.trans_up_1_12\
        );

    \I__621\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3538\,
            I => \d1.trans_up_1_9\
        );

    \I__619\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3532\,
            I => \d1.trans_up_sx\
        );

    \I__617\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3517\
        );

    \I__616\ : InMux
    port map (
            O => \N__3528\,
            I => \N__3517\
        );

    \I__615\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3517\
        );

    \I__614\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3517\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3517\,
            I => \d1.stateZ0\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__3514\,
            I => \N__3510\
        );

    \I__611\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3507\
        );

    \I__610\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3504\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3507\,
            I => \d1.syncZ0Z_1\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3504\,
            I => \d1.syncZ0Z_1\
        );

    \I__607\ : IoInMux
    port map (
            O => \N__3499\,
            I => \N__3496\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__605\ : Span12Mux_s8_h
    port map (
            O => \N__3493\,
            I => \N__3490\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__3490\,
            I => \d1.idle_i\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__602\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3481\,
            I => \state_RNIU5D07\
        );

    \I__600\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3475\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3475\,
            I => \state_RNIPC4P3_1\
        );

    \I__598\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3469\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3469\,
            I => \state_RNIPC4P3_8\
        );

    \I__596\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3448\
        );

    \I__595\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3448\
        );

    \I__594\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3448\
        );

    \I__593\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3441\
        );

    \I__592\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3441\
        );

    \I__591\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3441\
        );

    \I__590\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3438\
        );

    \I__589\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3431\
        );

    \I__588\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3431\
        );

    \I__587\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3431\
        );

    \I__586\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3426\
        );

    \I__585\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3426\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3448\,
            I => d2_trans_up_1
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3441\,
            I => d2_trans_up_1
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3438\,
            I => d2_trans_up_1
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3431\,
            I => d2_trans_up_1
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3426\,
            I => d2_trans_up_1
        );

    \I__579\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3412\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3412\,
            I => \state_RNIPC4P3_5\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3409\,
            I => \d1.count_RNI2PCEZ0Z_3_cascade_\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__3406\,
            I => \d1.trans_up_1_14_cascade_\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \N__3400\
        );

    \I__574\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3391\
        );

    \I__573\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3391\
        );

    \I__572\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3391\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3391\,
            I => s_up
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__3388\,
            I => \s_up_cascade_\
        );

    \I__569\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3378\
        );

    \I__568\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3378\
        );

    \I__567\ : InMux
    port map (
            O => \N__3383\,
            I => \N__3375\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3378\,
            I => s_dn_i
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3375\,
            I => s_dn_i
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__563\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3364\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3364\,
            I => \state_RNIU5D07_0\
        );

    \I__561\ : InMux
    port map (
            O => \N__3361\,
            I => \N__3358\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3358\,
            I => \state_RNIPC4P3_0\
        );

    \I__559\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3352\,
            I => \state_RNIPC4P3_2\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3349\,
            I => \d2.trans_up_1_12_cascade_\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__3346\,
            I => \d2.trans_up_1_sx_cascade_\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3343\,
            I => \d2_trans_up_1_cascade_\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__553\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3332\
        );

    \I__552\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3326\
        );

    \I__551\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3326\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3332\,
            I => \N__3323\
        );

    \I__549\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3320\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3315\
        );

    \I__547\ : Span4Mux_h
    port map (
            O => \N__3323\,
            I => \N__3315\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3320\,
            I => \pulse_lenZ0Z_2\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__3315\,
            I => \pulse_lenZ0Z_2\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3310\,
            I => \s_dn_i_cascade_\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3307\,
            I => \N__3304\
        );

    \I__542\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3301\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3301\,
            I => \un1_pulse_len_cry_2_c_RNOZ0\
        );

    \I__540\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3295\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3295\,
            I => \state_RNIPC4P3_3\
        );

    \I__538\ : InMux
    port map (
            O => \N__3292\,
            I => \p.count_1_cry_7\
        );

    \I__537\ : InMux
    port map (
            O => \N__3289\,
            I => \bfn_7_13_0_\
        );

    \I__536\ : InMux
    port map (
            O => \N__3286\,
            I => \p.count_1_cry_9\
        );

    \I__535\ : InMux
    port map (
            O => \N__3283\,
            I => \p.count_1_cry_10\
        );

    \I__534\ : InMux
    port map (
            O => \N__3280\,
            I => \p.count_1_cry_11\
        );

    \I__533\ : InMux
    port map (
            O => \N__3277\,
            I => \p.count_1_cry_12\
        );

    \I__532\ : InMux
    port map (
            O => \N__3274\,
            I => \p.count_1_cry_13\
        );

    \I__531\ : InMux
    port map (
            O => \N__3271\,
            I => \p.count_1_cry_14\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__529\ : InMux
    port map (
            O => \N__3265\,
            I => \N__3261\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__3264\,
            I => \N__3258\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3261\,
            I => \N__3255\
        );

    \I__526\ : InMux
    port map (
            O => \N__3258\,
            I => \N__3252\
        );

    \I__525\ : Span4Mux_h
    port map (
            O => \N__3255\,
            I => \N__3249\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3252\,
            I => \pulse_lenZ0Z_15\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__3249\,
            I => \pulse_lenZ0Z_15\
        );

    \I__522\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3241\,
            I => \p.count_i_15\
        );

    \I__520\ : InMux
    port map (
            O => \N__3238\,
            I => \p.CONTROL_PIN_2\
        );

    \I__519\ : IoInMux
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__517\ : IoSpan4Mux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__516\ : Sp12to4
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__515\ : Span12Mux_h
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__514\ : Span12Mux_v
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__3217\,
            I => \CONTROL_PIN_c\
        );

    \I__512\ : InMux
    port map (
            O => \N__3214\,
            I => \p.count_1_cry_1\
        );

    \I__511\ : InMux
    port map (
            O => \N__3211\,
            I => \p.count_1_cry_2\
        );

    \I__510\ : InMux
    port map (
            O => \N__3208\,
            I => \p.count_1_cry_3\
        );

    \I__509\ : InMux
    port map (
            O => \N__3205\,
            I => \p.count_1_cry_4\
        );

    \I__508\ : InMux
    port map (
            O => \N__3202\,
            I => \p.count_1_cry_5\
        );

    \I__507\ : InMux
    port map (
            O => \N__3199\,
            I => \p.count_1_cry_6\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__3196\,
            I => \N__3193\
        );

    \I__505\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3189\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3192\,
            I => \N__3186\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3189\,
            I => \N__3183\
        );

    \I__502\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__501\ : Span4Mux_h
    port map (
            O => \N__3183\,
            I => \N__3177\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3180\,
            I => \pulse_lenZ0Z_7\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__3177\,
            I => \pulse_lenZ0Z_7\
        );

    \I__498\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3169\,
            I => \p.count_i_7\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3166\,
            I => \N__3162\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__3165\,
            I => \N__3159\
        );

    \I__494\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3156\
        );

    \I__493\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3153\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3156\,
            I => \N__3150\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3153\,
            I => \N__3145\
        );

    \I__490\ : Span4Mux_h
    port map (
            O => \N__3150\,
            I => \N__3145\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__3145\,
            I => \pulse_lenZ0Z_8\
        );

    \I__488\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3139\,
            I => \p.count_i_8\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__3136\,
            I => \N__3132\
        );

    \I__485\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3129\
        );

    \I__484\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3126\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3129\,
            I => \N__3123\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3126\,
            I => \pulse_lenZ0Z_9\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3123\,
            I => \pulse_lenZ0Z_9\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3118\,
            I => \N__3115\
        );

    \I__479\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3112\,
            I => \p.count_i_9\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__3109\,
            I => \N__3105\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__3108\,
            I => \N__3102\
        );

    \I__475\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3099\
        );

    \I__474\ : InMux
    port map (
            O => \N__3102\,
            I => \N__3096\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3099\,
            I => \N__3093\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3096\,
            I => \pulse_lenZ0Z_10\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3093\,
            I => \pulse_lenZ0Z_10\
        );

    \I__470\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3085\,
            I => \p.count_i_10\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__467\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3075\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3078\,
            I => \N__3072\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3075\,
            I => \N__3069\
        );

    \I__464\ : InMux
    port map (
            O => \N__3072\,
            I => \N__3066\
        );

    \I__463\ : Span4Mux_h
    port map (
            O => \N__3069\,
            I => \N__3063\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3066\,
            I => \pulse_lenZ0Z_11\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__3063\,
            I => \pulse_lenZ0Z_11\
        );

    \I__460\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3055\,
            I => \p.count_i_11\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3052\,
            I => \N__3048\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3051\,
            I => \N__3045\
        );

    \I__456\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3042\
        );

    \I__455\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3039\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3042\,
            I => \N__3036\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3039\,
            I => \pulse_lenZ0Z_12\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__3036\,
            I => \pulse_lenZ0Z_12\
        );

    \I__451\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3028\,
            I => \p.count_i_12\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__3025\,
            I => \N__3021\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__3024\,
            I => \N__3018\
        );

    \I__447\ : InMux
    port map (
            O => \N__3021\,
            I => \N__3015\
        );

    \I__446\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3012\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3015\,
            I => \N__3009\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3012\,
            I => \pulse_lenZ0Z_13\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__3009\,
            I => \pulse_lenZ0Z_13\
        );

    \I__442\ : InMux
    port map (
            O => \N__3004\,
            I => \N__3001\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3001\,
            I => \p.count_i_13\
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__2998\,
            I => \N__2994\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__2997\,
            I => \N__2991\
        );

    \I__438\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2988\
        );

    \I__437\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2985\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2982\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2985\,
            I => \pulse_lenZ0Z_14\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__2982\,
            I => \pulse_lenZ0Z_14\
        );

    \I__433\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2974\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2974\,
            I => \p.count_i_14\
        );

    \I__431\ : InMux
    port map (
            O => \N__2971\,
            I => un1_pulse_len_cry_14
        );

    \I__430\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2965\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2965\,
            I => \state_RNIPC4P3_4\
        );

    \I__428\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2959\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2959\,
            I => \state_RNIPC4P3_7\
        );

    \I__426\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2953\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2953\,
            I => \p.count_i_2\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__2950\,
            I => \N__2947\
        );

    \I__423\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2943\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__2946\,
            I => \N__2940\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2943\,
            I => \N__2937\
        );

    \I__420\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2934\
        );

    \I__419\ : Span4Mux_h
    port map (
            O => \N__2937\,
            I => \N__2931\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2934\,
            I => \pulse_lenZ0Z_3\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__2931\,
            I => \pulse_lenZ0Z_3\
        );

    \I__416\ : InMux
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2923\,
            I => \p.count_i_3\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2920\,
            I => \N__2916\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2919\,
            I => \N__2913\
        );

    \I__412\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2910\
        );

    \I__411\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2907\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2910\,
            I => \N__2904\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2907\,
            I => \pulse_lenZ0Z_4\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__2904\,
            I => \pulse_lenZ0Z_4\
        );

    \I__407\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2896\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2896\,
            I => \p.count_i_4\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__2893\,
            I => \N__2890\
        );

    \I__404\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2887\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2887\,
            I => \N__2883\
        );

    \I__402\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2880\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__2883\,
            I => \N__2877\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2880\,
            I => \pulse_lenZ0Z_5\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__2877\,
            I => \pulse_lenZ0Z_5\
        );

    \I__398\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2869\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2869\,
            I => \p.count_i_5\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__2866\,
            I => \N__2863\
        );

    \I__395\ : InMux
    port map (
            O => \N__2863\,
            I => \N__2859\
        );

    \I__394\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2856\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2859\,
            I => \N__2853\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2856\,
            I => \pulse_lenZ0Z_6\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__2853\,
            I => \pulse_lenZ0Z_6\
        );

    \I__390\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2845\,
            I => \p.count_i_6\
        );

    \I__388\ : InMux
    port map (
            O => \N__2842\,
            I => un1_pulse_len_cry_5
        );

    \I__387\ : InMux
    port map (
            O => \N__2839\,
            I => un1_pulse_len_cry_6
        );

    \I__386\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2833\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2833\,
            I => \state_RNIPC4P3_6\
        );

    \I__384\ : InMux
    port map (
            O => \N__2830\,
            I => un1_pulse_len_cry_7
        );

    \I__383\ : InMux
    port map (
            O => \N__2827\,
            I => un1_pulse_len_cry_8
        );

    \I__382\ : InMux
    port map (
            O => \N__2824\,
            I => \bfn_7_9_0_\
        );

    \I__381\ : InMux
    port map (
            O => \N__2821\,
            I => un1_pulse_len_cry_10
        );

    \I__380\ : InMux
    port map (
            O => \N__2818\,
            I => un1_pulse_len_cry_11
        );

    \I__379\ : InMux
    port map (
            O => \N__2815\,
            I => un1_pulse_len_cry_12
        );

    \I__378\ : InMux
    port map (
            O => \N__2812\,
            I => un1_pulse_len_cry_13
        );

    \I__377\ : InMux
    port map (
            O => \N__2809\,
            I => \N__2806\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2806\,
            I => \p.prescaler_1_cry_5_THRU_CO\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__2803\,
            I => \N__2798\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__2802\,
            I => \N__2795\
        );

    \I__373\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2792\
        );

    \I__372\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2787\
        );

    \I__371\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2787\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2792\,
            I => \p.prescalerZ0Z_6\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2787\,
            I => \p.prescalerZ0Z_6\
        );

    \I__368\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2779\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2779\,
            I => \p.prescaler_1_cry_4_THRU_CO\
        );

    \I__366\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2771\
        );

    \I__365\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2766\
        );

    \I__364\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2766\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2771\,
            I => \p.prescalerZ0Z_5\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2766\,
            I => \p.prescalerZ0Z_5\
        );

    \I__361\ : InMux
    port map (
            O => \N__2761\,
            I => \N__2755\
        );

    \I__360\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2748\
        );

    \I__359\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2748\
        );

    \I__358\ : InMux
    port map (
            O => \N__2758\,
            I => \N__2748\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2755\,
            I => \p.prescalerZ0Z_0\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2748\,
            I => \p.prescalerZ0Z_0\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__354\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2735\
        );

    \I__353\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2730\
        );

    \I__352\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2730\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2735\,
            I => \p.prescalerZ0Z_1\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2730\,
            I => \p.prescalerZ0Z_1\
        );

    \I__349\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2722\,
            I => \state_RNIPC4P3\
        );

    \I__347\ : InMux
    port map (
            O => \N__2719\,
            I => un1_pulse_len_cry_2
        );

    \I__346\ : InMux
    port map (
            O => \N__2716\,
            I => un1_pulse_len_cry_3
        );

    \I__345\ : InMux
    port map (
            O => \N__2713\,
            I => un1_pulse_len_cry_4
        );

    \I__344\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2706\
        );

    \I__343\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2703\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2706\,
            I => \p.prescalerZ0Z_20\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2703\,
            I => \p.prescalerZ0Z_20\
        );

    \I__340\ : InMux
    port map (
            O => \N__2698\,
            I => \p.prescaler_1_cry_19\
        );

    \I__339\ : InMux
    port map (
            O => \N__2695\,
            I => \N__2691\
        );

    \I__338\ : InMux
    port map (
            O => \N__2694\,
            I => \N__2688\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2691\,
            I => \p.prescalerZ0Z_21\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2688\,
            I => \p.prescalerZ0Z_21\
        );

    \I__335\ : InMux
    port map (
            O => \N__2683\,
            I => \p.prescaler_1_cry_20\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__2680\,
            I => \N__2676\
        );

    \I__333\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2673\
        );

    \I__332\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2670\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2673\,
            I => \p.prescalerZ0Z_22\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2670\,
            I => \p.prescalerZ0Z_22\
        );

    \I__329\ : InMux
    port map (
            O => \N__2665\,
            I => \p.prescaler_1_cry_21\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2662\,
            I => \N__2658\
        );

    \I__327\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2655\
        );

    \I__326\ : InMux
    port map (
            O => \N__2658\,
            I => \N__2652\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2655\,
            I => \p.prescalerZ0Z_23\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2652\,
            I => \p.prescalerZ0Z_23\
        );

    \I__323\ : InMux
    port map (
            O => \N__2647\,
            I => \p.prescaler_1_cry_22\
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__2644\,
            I => \N__2641\
        );

    \I__321\ : InMux
    port map (
            O => \N__2641\,
            I => \N__2637\
        );

    \I__320\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2634\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2637\,
            I => \N__2631\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2634\,
            I => \p.prescalerZ0Z_24\
        );

    \I__317\ : Odrv4
    port map (
            O => \N__2631\,
            I => \p.prescalerZ0Z_24\
        );

    \I__316\ : InMux
    port map (
            O => \N__2626\,
            I => \p.prescaler_1_cry_23\
        );

    \I__315\ : CascadeMux
    port map (
            O => \N__2623\,
            I => \N__2620\
        );

    \I__314\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2616\
        );

    \I__313\ : InMux
    port map (
            O => \N__2619\,
            I => \N__2613\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2616\,
            I => \N__2610\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2613\,
            I => \p.prescalerZ0Z_25\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__2610\,
            I => \p.prescalerZ0Z_25\
        );

    \I__309\ : InMux
    port map (
            O => \N__2605\,
            I => \bfn_2_14_0_\
        );

    \I__308\ : InMux
    port map (
            O => \N__2602\,
            I => \p.prescaler_1_cry_25\
        );

    \I__307\ : CascadeMux
    port map (
            O => \N__2599\,
            I => \N__2595\
        );

    \I__306\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2592\
        );

    \I__305\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2589\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2592\,
            I => \p.prescalerZ0Z_26\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2589\,
            I => \p.prescalerZ0Z_26\
        );

    \I__302\ : InMux
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2581\,
            I => \N__2578\
        );

    \I__300\ : Odrv4
    port map (
            O => \N__2578\,
            I => \p.prescaler12_0_and\
        );

    \I__299\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2571\
        );

    \I__298\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2568\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2571\,
            I => \p.prescalerZ0Z_12\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2568\,
            I => \p.prescalerZ0Z_12\
        );

    \I__295\ : InMux
    port map (
            O => \N__2563\,
            I => \p.prescaler_1_cry_11\
        );

    \I__294\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2556\
        );

    \I__293\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2553\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2556\,
            I => \p.prescalerZ0Z_13\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2553\,
            I => \p.prescalerZ0Z_13\
        );

    \I__290\ : InMux
    port map (
            O => \N__2548\,
            I => \p.prescaler_1_cry_12\
        );

    \I__289\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2541\
        );

    \I__288\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2538\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2541\,
            I => \p.prescalerZ0Z_14\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2538\,
            I => \p.prescalerZ0Z_14\
        );

    \I__285\ : InMux
    port map (
            O => \N__2533\,
            I => \p.prescaler_1_cry_13\
        );

    \I__284\ : InMux
    port map (
            O => \N__2530\,
            I => \N__2526\
        );

    \I__283\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2523\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2526\,
            I => \p.prescalerZ0Z_15\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2523\,
            I => \p.prescalerZ0Z_15\
        );

    \I__280\ : InMux
    port map (
            O => \N__2518\,
            I => \p.prescaler_1_cry_14\
        );

    \I__279\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2511\
        );

    \I__278\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2508\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2511\,
            I => \p.prescalerZ0Z_16\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2508\,
            I => \p.prescalerZ0Z_16\
        );

    \I__275\ : InMux
    port map (
            O => \N__2503\,
            I => \p.prescaler_1_cry_15\
        );

    \I__274\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2496\
        );

    \I__273\ : InMux
    port map (
            O => \N__2499\,
            I => \N__2493\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2496\,
            I => \p.prescalerZ0Z_17\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2493\,
            I => \p.prescalerZ0Z_17\
        );

    \I__270\ : InMux
    port map (
            O => \N__2488\,
            I => \bfn_2_13_0_\
        );

    \I__269\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2481\
        );

    \I__268\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2478\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2481\,
            I => \N__2475\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2478\,
            I => \p.prescalerZ0Z_18\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2475\,
            I => \p.prescalerZ0Z_18\
        );

    \I__264\ : InMux
    port map (
            O => \N__2470\,
            I => \p.prescaler_1_cry_17\
        );

    \I__263\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2463\
        );

    \I__262\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2460\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2463\,
            I => \p.prescalerZ0Z_19\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2460\,
            I => \p.prescalerZ0Z_19\
        );

    \I__259\ : InMux
    port map (
            O => \N__2455\,
            I => \p.prescaler_1_cry_18\
        );

    \I__258\ : InMux
    port map (
            O => \N__2452\,
            I => \N__2448\
        );

    \I__257\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2445\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2448\,
            I => \p.prescalerZ0Z_3\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2445\,
            I => \p.prescalerZ0Z_3\
        );

    \I__254\ : InMux
    port map (
            O => \N__2440\,
            I => \p.prescaler_1_cry_2\
        );

    \I__253\ : InMux
    port map (
            O => \N__2437\,
            I => \N__2433\
        );

    \I__252\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2430\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2433\,
            I => \p.prescalerZ0Z_4\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2430\,
            I => \p.prescalerZ0Z_4\
        );

    \I__249\ : InMux
    port map (
            O => \N__2425\,
            I => \p.prescaler_1_cry_3\
        );

    \I__248\ : InMux
    port map (
            O => \N__2422\,
            I => \p.prescaler_1_cry_4\
        );

    \I__247\ : InMux
    port map (
            O => \N__2419\,
            I => \p.prescaler_1_cry_5\
        );

    \I__246\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2412\
        );

    \I__245\ : InMux
    port map (
            O => \N__2415\,
            I => \N__2409\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2412\,
            I => \p.prescalerZ0Z_7\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2409\,
            I => \p.prescalerZ0Z_7\
        );

    \I__242\ : InMux
    port map (
            O => \N__2404\,
            I => \p.prescaler_1_cry_6\
        );

    \I__241\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2397\
        );

    \I__240\ : InMux
    port map (
            O => \N__2400\,
            I => \N__2394\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2397\,
            I => \p.prescalerZ0Z_8\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2394\,
            I => \p.prescalerZ0Z_8\
        );

    \I__237\ : InMux
    port map (
            O => \N__2389\,
            I => \p.prescaler_1_cry_7\
        );

    \I__236\ : InMux
    port map (
            O => \N__2386\,
            I => \N__2382\
        );

    \I__235\ : InMux
    port map (
            O => \N__2385\,
            I => \N__2379\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2382\,
            I => \p.prescalerZ0Z_9\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2379\,
            I => \p.prescalerZ0Z_9\
        );

    \I__232\ : InMux
    port map (
            O => \N__2374\,
            I => \bfn_2_12_0_\
        );

    \I__231\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2367\
        );

    \I__230\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2364\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2367\,
            I => \p.prescalerZ0Z_10\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2364\,
            I => \p.prescalerZ0Z_10\
        );

    \I__227\ : InMux
    port map (
            O => \N__2359\,
            I => \p.prescaler_1_cry_9\
        );

    \I__226\ : InMux
    port map (
            O => \N__2356\,
            I => \N__2352\
        );

    \I__225\ : InMux
    port map (
            O => \N__2355\,
            I => \N__2349\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2352\,
            I => \p.prescalerZ0Z_11\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2349\,
            I => \p.prescalerZ0Z_11\
        );

    \I__222\ : InMux
    port map (
            O => \N__2344\,
            I => \p.prescaler_1_cry_10\
        );

    \I__221\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2338\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2338\,
            I => \p.prescaler12_4_and\
        );

    \I__219\ : InMux
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2332\,
            I => \p.prescaler12_2_and\
        );

    \I__217\ : InMux
    port map (
            O => \N__2329\,
            I => \N__2326\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__2326\,
            I => \p.prescaler12_6_and\
        );

    \I__215\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2320\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2320\,
            I => \p.prescaler12_5_and\
        );

    \I__213\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2314\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2314\,
            I => \p.prescaler12_3_and\
        );

    \I__211\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2308\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2308\,
            I => \N__2305\
        );

    \I__209\ : Odrv4
    port map (
            O => \N__2305\,
            I => \p.prescaler12_1_and\
        );

    \I__208\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2297\
        );

    \I__207\ : InMux
    port map (
            O => \N__2301\,
            I => \N__2292\
        );

    \I__206\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2292\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2297\,
            I => \p.prescalerZ0Z_2\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2292\,
            I => \p.prescalerZ0Z_2\
        );

    \I__203\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2284\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__2284\,
            I => \p.prescaler_1_cry_1_THRU_CO\
        );

    \I__201\ : InMux
    port map (
            O => \N__2281\,
            I => \p.prescaler_1_cry_1\
        );

    \I__200\ : InMux
    port map (
            O => \N__2278\,
            I => \p.prescaler12\
        );

    \I__199\ : IoInMux
    port map (
            O => \N__2275\,
            I => \N__2272\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__2272\,
            I => \N__2269\
        );

    \I__197\ : Odrv12
    port map (
            O => \N__2269\,
            I => \p.prescaler12_THRU_CO\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_pulse_len_cry_9,
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \p.prescaler_1_cry_8\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \p.prescaler_1_cry_16\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \p.prescaler_1_cry_24\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \p.count_1_cry_8\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d2.un3_count_cry_8\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \d1.un3_count_cry_8\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \p.CONTROL_PIN_2_cry_9\,
            carryinitout => \bfn_7_11_0_\
        );

    \p.prescaler12_6_c_RNIPKT\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2275\,
            GLOBALBUFFEROUTPUT => \p.prescaler12_g\
        );

    \d2.sync_1_RNIMV5K_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4030\,
            GLOBALBUFFEROUTPUT => \d2.idle_i_g\
        );

    \d1.sync_1_RNIKI1C_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3499\,
            GLOBALBUFFEROUTPUT => \d1.idle_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \p.prescaler12_0_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2584\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \p.prescaler12_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_1_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2311\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_0\,
            carryout => \p.prescaler12_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_2_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2335\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_1\,
            carryout => \p.prescaler12_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_3_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2317\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_2\,
            carryout => \p.prescaler12_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_4_c_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2341\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_3\,
            carryout => \p.prescaler12_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_5_c_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2323\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_4\,
            carryout => \p.prescaler12_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_6_c_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \p.prescaler12_5\,
            carryout => \p.prescaler12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_THRU_LUT4_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2278\,
            lcout => \p.prescaler12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_4_c_RNO_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2385\,
            in1 => \N__2355\,
            in2 => \N__2680\,
            in3 => \N__2451\,
            lcout => \p.prescaler12_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2287\,
            in1 => \N__2301\,
            in2 => \_gnd_net_\,
            in3 => \N__4439\,
            lcout => \p.prescalerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_2_c_RNO_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2499\,
            in1 => \N__2559\,
            in2 => \N__2623\,
            in3 => \N__2574\,
            lcout => \p.prescaler12_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_6_c_RNO_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2466\,
            in1 => \N__2514\,
            in2 => \_gnd_net_\,
            in3 => \N__2415\,
            lcout => \p.prescaler12_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_5_c_RNO_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2529\,
            in1 => \N__2400\,
            in2 => \N__2644\,
            in3 => \N__2436\,
            lcout => \p.prescaler12_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_3_c_RNO_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2370\,
            in1 => \N__2485\,
            in2 => \N__2662\,
            in3 => \N__2300\,
            lcout => \p.prescaler12_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_1_c_RNO_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2694\,
            in1 => \N__2709\,
            in2 => \N__2599\,
            in3 => \N__2544\,
            lcout => \p.prescaler12_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_1_cry_1_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2761\,
            in2 => \N__2743\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \p.prescaler_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_1_cry_1_THRU_LUT4_0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2302\,
            in2 => \_gnd_net_\,
            in3 => \N__2281\,
            lcout => \p.prescaler_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_1\,
            carryout => \p.prescaler_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_3_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2452\,
            in2 => \_gnd_net_\,
            in3 => \N__2440\,
            lcout => \p.prescalerZ0Z_3\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_2\,
            carryout => \p.prescaler_1_cry_3\,
            clk => \N__4813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_4_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2437\,
            in2 => \_gnd_net_\,
            in3 => \N__2425\,
            lcout => \p.prescalerZ0Z_4\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_3\,
            carryout => \p.prescaler_1_cry_4\,
            clk => \N__4813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_1_cry_4_THRU_LUT4_0_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2776\,
            in2 => \_gnd_net_\,
            in3 => \N__2422\,
            lcout => \p.prescaler_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_4\,
            carryout => \p.prescaler_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_1_cry_5_THRU_LUT4_0_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2801\,
            in2 => \_gnd_net_\,
            in3 => \N__2419\,
            lcout => \p.prescaler_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_5\,
            carryout => \p.prescaler_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_7_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2416\,
            in2 => \_gnd_net_\,
            in3 => \N__2404\,
            lcout => \p.prescalerZ0Z_7\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_6\,
            carryout => \p.prescaler_1_cry_7\,
            clk => \N__4813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2401\,
            in2 => \_gnd_net_\,
            in3 => \N__2389\,
            lcout => \p.prescalerZ0Z_8\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_7\,
            carryout => \p.prescaler_1_cry_8\,
            clk => \N__4813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_9_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2386\,
            in2 => \_gnd_net_\,
            in3 => \N__2374\,
            lcout => \p.prescalerZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \p.prescaler_1_cry_9\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_10_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2371\,
            in2 => \_gnd_net_\,
            in3 => \N__2359\,
            lcout => \p.prescalerZ0Z_10\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_9\,
            carryout => \p.prescaler_1_cry_10\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_11_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2356\,
            in2 => \_gnd_net_\,
            in3 => \N__2344\,
            lcout => \p.prescalerZ0Z_11\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_10\,
            carryout => \p.prescaler_1_cry_11\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_12_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2575\,
            in2 => \_gnd_net_\,
            in3 => \N__2563\,
            lcout => \p.prescalerZ0Z_12\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_11\,
            carryout => \p.prescaler_1_cry_12\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_13_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2560\,
            in2 => \_gnd_net_\,
            in3 => \N__2548\,
            lcout => \p.prescalerZ0Z_13\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_12\,
            carryout => \p.prescaler_1_cry_13\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_14_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2545\,
            in2 => \_gnd_net_\,
            in3 => \N__2533\,
            lcout => \p.prescalerZ0Z_14\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_13\,
            carryout => \p.prescaler_1_cry_14\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_15_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2530\,
            in2 => \_gnd_net_\,
            in3 => \N__2518\,
            lcout => \p.prescalerZ0Z_15\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_14\,
            carryout => \p.prescaler_1_cry_15\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_16_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2515\,
            in2 => \_gnd_net_\,
            in3 => \N__2503\,
            lcout => \p.prescalerZ0Z_16\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_15\,
            carryout => \p.prescaler_1_cry_16\,
            clk => \N__4809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_17_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2500\,
            in2 => \_gnd_net_\,
            in3 => \N__2488\,
            lcout => \p.prescalerZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \p.prescaler_1_cry_17\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_18_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2484\,
            in2 => \_gnd_net_\,
            in3 => \N__2470\,
            lcout => \p.prescalerZ0Z_18\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_17\,
            carryout => \p.prescaler_1_cry_18\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_19_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2467\,
            in2 => \_gnd_net_\,
            in3 => \N__2455\,
            lcout => \p.prescalerZ0Z_19\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_18\,
            carryout => \p.prescaler_1_cry_19\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_20_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2710\,
            in2 => \_gnd_net_\,
            in3 => \N__2698\,
            lcout => \p.prescalerZ0Z_20\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_19\,
            carryout => \p.prescaler_1_cry_20\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_21_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2695\,
            in2 => \_gnd_net_\,
            in3 => \N__2683\,
            lcout => \p.prescalerZ0Z_21\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_20\,
            carryout => \p.prescaler_1_cry_21\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_22_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2679\,
            in2 => \_gnd_net_\,
            in3 => \N__2665\,
            lcout => \p.prescalerZ0Z_22\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_21\,
            carryout => \p.prescaler_1_cry_22\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_23_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2661\,
            in2 => \_gnd_net_\,
            in3 => \N__2647\,
            lcout => \p.prescalerZ0Z_23\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_22\,
            carryout => \p.prescaler_1_cry_23\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_24_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2640\,
            in2 => \_gnd_net_\,
            in3 => \N__2626\,
            lcout => \p.prescalerZ0Z_24\,
            ltout => OPEN,
            carryin => \p.prescaler_1_cry_23\,
            carryout => \p.prescaler_1_cry_24\,
            clk => \N__4808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_25_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2619\,
            in2 => \_gnd_net_\,
            in3 => \N__2605\,
            lcout => \p.prescalerZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \p.prescaler_1_cry_25\,
            clk => \N__4805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_26_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2598\,
            in2 => \_gnd_net_\,
            in3 => \N__2602\,
            lcout => \p.prescalerZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_0_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \p.prescalerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler12_0_c_RNO_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2774\,
            in1 => \N__2738\,
            in2 => \N__2802\,
            in3 => \N__2758\,
            lcout => \p.prescaler12_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_6_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__4441\,
            in1 => \_gnd_net_\,
            in2 => \N__2803\,
            in3 => \N__2809\,
            lcout => \p.prescalerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_5_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2782\,
            in1 => \N__2775\,
            in2 => \_gnd_net_\,
            in3 => \N__4440\,
            lcout => \p.prescalerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.prescaler_1_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2739\,
            in2 => \_gnd_net_\,
            in3 => \N__2760\,
            lcout => \p.prescalerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4084\,
            lcout => \state_RNIPC4P3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4076\,
            in2 => \_gnd_net_\,
            in3 => \N__3455\,
            lcout => \state_RNIPC4P3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_pulse_len_cry_2_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3331\,
            in2 => \N__3307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => un1_pulse_len_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2725\,
            in2 => \N__2946\,
            in3 => \N__2719\,
            lcout => \pulse_lenZ0Z_3\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_2,
            carryout => un1_pulse_len_cry_3,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_4_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3361\,
            in2 => \N__2919\,
            in3 => \N__2716\,
            lcout => \pulse_lenZ0Z_4\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_3,
            carryout => un1_pulse_len_cry_4,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2886\,
            in2 => \N__3370\,
            in3 => \N__2713\,
            lcout => \pulse_lenZ0Z_5\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_4,
            carryout => un1_pulse_len_cry_5,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_6_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2862\,
            in2 => \N__3487\,
            in3 => \N__2842\,
            lcout => \pulse_lenZ0Z_6\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_5,
            carryout => un1_pulse_len_cry_6,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_7_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3298\,
            in2 => \N__3192\,
            in3 => \N__2839\,
            lcout => \pulse_lenZ0Z_7\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_6,
            carryout => un1_pulse_len_cry_7,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_8_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2836\,
            in2 => \N__3165\,
            in3 => \N__2830\,
            lcout => \pulse_lenZ0Z_8\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_7,
            carryout => un1_pulse_len_cry_8,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_9_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3355\,
            in2 => \N__3136\,
            in3 => \N__2827\,
            lcout => \pulse_lenZ0Z_9\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_8,
            carryout => un1_pulse_len_cry_9,
            clk => \N__4806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_10_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3478\,
            in2 => \N__3108\,
            in3 => \N__2824\,
            lcout => \pulse_lenZ0Z_10\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => un1_pulse_len_cry_10,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_11_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3415\,
            in2 => \N__3078\,
            in3 => \N__2821\,
            lcout => \pulse_lenZ0Z_11\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_10,
            carryout => un1_pulse_len_cry_11,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_12_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2962\,
            in2 => \N__3051\,
            in3 => \N__2818\,
            lcout => \pulse_lenZ0Z_12\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_11,
            carryout => un1_pulse_len_cry_12,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_13_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2968\,
            in2 => \N__3024\,
            in3 => \N__2815\,
            lcout => \pulse_lenZ0Z_13\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_12,
            carryout => un1_pulse_len_cry_13,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_14_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3472\,
            in2 => \N__2997\,
            in3 => \N__2812\,
            lcout => \pulse_lenZ0Z_14\,
            ltout => OPEN,
            carryin => un1_pulse_len_cry_13,
            carryout => un1_pulse_len_cry_14,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_15_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__3466\,
            in2 => \N__3264\,
            in3 => \N__2971\,
            lcout => \pulse_lenZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_4_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3465\,
            in1 => \_gnd_net_\,
            in2 => \N__4116\,
            in3 => \_gnd_net_\,
            lcout => \state_RNIPC4P3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4108\,
            in2 => \_gnd_net_\,
            in3 => \N__3464\,
            lcout => \state_RNIPC4P3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_2_c_inv_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2956\,
            in2 => \N__3340\,
            in3 => \N__3622\,
            lcout => \p.count_i_2\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \p.CONTROL_PIN_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_3_c_inv_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2926\,
            in2 => \N__2950\,
            in3 => \N__3643\,
            lcout => \p.count_i_3\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_2\,
            carryout => \p.CONTROL_PIN_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_4_c_inv_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2899\,
            in2 => \N__2920\,
            in3 => \N__3703\,
            lcout => \p.count_i_4\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_3\,
            carryout => \p.CONTROL_PIN_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_5_c_inv_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2872\,
            in2 => \N__2893\,
            in3 => \N__3790\,
            lcout => \p.count_i_5\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_4\,
            carryout => \p.CONTROL_PIN_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_6_c_inv_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2848\,
            in2 => \N__2866\,
            in3 => \N__3877\,
            lcout => \p.count_i_6\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_5\,
            carryout => \p.CONTROL_PIN_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_7_c_inv_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3835\,
            in1 => \N__3172\,
            in2 => \N__3196\,
            in3 => \_gnd_net_\,
            lcout => \p.count_i_7\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_6\,
            carryout => \p.CONTROL_PIN_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_8_c_inv_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3142\,
            in2 => \N__3166\,
            in3 => \N__3922\,
            lcout => \p.count_i_8\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_7\,
            carryout => \p.CONTROL_PIN_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_9_c_inv_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3135\,
            in2 => \N__3118\,
            in3 => \N__3748\,
            lcout => \p.count_i_9\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_8\,
            carryout => \p.CONTROL_PIN_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_10_c_inv_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3088\,
            in2 => \N__3109\,
            in3 => \N__3769\,
            lcout => \p.count_i_10\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \p.CONTROL_PIN_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_11_c_inv_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3058\,
            in2 => \N__3082\,
            in3 => \N__3726\,
            lcout => \p.count_i_11\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_10\,
            carryout => \p.CONTROL_PIN_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_12_c_inv_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3031\,
            in2 => \N__3052\,
            in3 => \N__3856\,
            lcout => \p.count_i_12\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_11\,
            carryout => \p.CONTROL_PIN_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_13_c_inv_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3004\,
            in2 => \N__3025\,
            in3 => \N__3813\,
            lcout => \p.count_i_13\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_12\,
            carryout => \p.CONTROL_PIN_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_14_c_inv_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2977\,
            in2 => \N__2998\,
            in3 => \N__3943\,
            lcout => \p.count_i_14\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_13\,
            carryout => \p.CONTROL_PIN_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_2_cry_15_c_inv_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3901\,
            in1 => \N__3244\,
            in2 => \N__3268\,
            in3 => \_gnd_net_\,
            lcout => \p.count_i_15\,
            ltout => OPEN,
            carryin => \p.CONTROL_PIN_2_cry_14\,
            carryout => \p.CONTROL_PIN_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.CONTROL_PIN_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3238\,
            lcout => \CONTROL_PIN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4797\,
            ce => \N__4427\,
            sr => \_gnd_net_\
        );

    \p.count_1_cry_1_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4465\,
            in2 => \N__4492\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \p.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.count_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3621\,
            in2 => \_gnd_net_\,
            in3 => \N__3214\,
            lcout => \p.countZ0Z_2\,
            ltout => OPEN,
            carryin => \p.count_1_cry_1\,
            carryout => \p.count_1_cry_2\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_3_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3642\,
            in2 => \_gnd_net_\,
            in3 => \N__3211\,
            lcout => \p.countZ0Z_3\,
            ltout => OPEN,
            carryin => \p.count_1_cry_2\,
            carryout => \p.count_1_cry_3\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3702\,
            in2 => \_gnd_net_\,
            in3 => \N__3208\,
            lcout => \p.countZ0Z_4\,
            ltout => OPEN,
            carryin => \p.count_1_cry_3\,
            carryout => \p.count_1_cry_4\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3665\,
            in1 => \N__3789\,
            in2 => \_gnd_net_\,
            in3 => \N__3205\,
            lcout => \p.countZ0Z_5\,
            ltout => OPEN,
            carryin => \p.count_1_cry_4\,
            carryout => \p.count_1_cry_5\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_6_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__3202\,
            lcout => \p.countZ0Z_6\,
            ltout => OPEN,
            carryin => \p.count_1_cry_5\,
            carryout => \p.count_1_cry_6\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_7_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3834\,
            in2 => \_gnd_net_\,
            in3 => \N__3199\,
            lcout => \p.countZ0Z_7\,
            ltout => OPEN,
            carryin => \p.count_1_cry_6\,
            carryout => \p.count_1_cry_7\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_8_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3921\,
            in2 => \_gnd_net_\,
            in3 => \N__3292\,
            lcout => \p.countZ0Z_8\,
            ltout => OPEN,
            carryin => \p.count_1_cry_7\,
            carryout => \p.count_1_cry_8\,
            clk => \N__4793\,
            ce => \N__4428\,
            sr => \_gnd_net_\
        );

    \p.count_9_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3664\,
            in1 => \N__3747\,
            in2 => \_gnd_net_\,
            in3 => \N__3289\,
            lcout => \p.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \p.count_1_cry_9\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_10_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3666\,
            in1 => \N__3768\,
            in2 => \_gnd_net_\,
            in3 => \N__3286\,
            lcout => \p.countZ0Z_10\,
            ltout => OPEN,
            carryin => \p.count_1_cry_9\,
            carryout => \p.count_1_cry_10\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_11_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3663\,
            in1 => \N__3725\,
            in2 => \_gnd_net_\,
            in3 => \N__3283\,
            lcout => \p.countZ0Z_11\,
            ltout => OPEN,
            carryin => \p.count_1_cry_10\,
            carryout => \p.count_1_cry_11\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_12_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3855\,
            in2 => \_gnd_net_\,
            in3 => \N__3280\,
            lcout => \p.countZ0Z_12\,
            ltout => OPEN,
            carryin => \p.count_1_cry_11\,
            carryout => \p.count_1_cry_12\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_13_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3812\,
            in2 => \_gnd_net_\,
            in3 => \N__3277\,
            lcout => \p.countZ0Z_13\,
            ltout => OPEN,
            carryin => \p.count_1_cry_12\,
            carryout => \p.count_1_cry_13\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_14_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3667\,
            in1 => \N__3942\,
            in2 => \_gnd_net_\,
            in3 => \N__3274\,
            lcout => \p.countZ0Z_14\,
            ltout => OPEN,
            carryin => \p.count_1_cry_13\,
            carryout => \p.count_1_cry_14\,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \p.count_15_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3899\,
            in2 => \_gnd_net_\,
            in3 => \N__3271\,
            lcout => \p.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4792\,
            ce => \N__4429\,
            sr => \_gnd_net_\
        );

    \d2.state_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__3459\,
            in1 => \_gnd_net_\,
            in2 => \N__4102\,
            in3 => \_gnd_net_\,
            lcout => d2_state,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4077\,
            in2 => \_gnd_net_\,
            in3 => \N__3457\,
            lcout => \state_RNIPC4P3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3458\,
            in1 => \_gnd_net_\,
            in2 => \N__4101\,
            in3 => \_gnd_net_\,
            lcout => \state_RNIPC4P3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_len_2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__3385\,
            in1 => \_gnd_net_\,
            in2 => \N__3403\,
            in3 => \N__3335\,
            lcout => \pulse_lenZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNINDU8_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4396\,
            in2 => \_gnd_net_\,
            in3 => \N__4174\,
            lcout => OPEN,
            ltout => \d2.trans_up_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_RNI3PR51_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101111111"
        )
    port map (
            in0 => \N__4128\,
            in1 => \N__4370\,
            in2 => \N__3349\,
            in3 => \N__4073\,
            lcout => OPEN,
            ltout => \d2.trans_up_1_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIK9TB3_10_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3595\,
            in1 => \N__3583\,
            in2 => \N__3346\,
            in3 => \N__4186\,
            lcout => d2_trans_up_1,
            ltout => \d2_trans_up_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_9_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3343\,
            in3 => \N__4074\,
            lcout => s_dn_i,
            ltout => \s_dn_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_pulse_len_cry_2_c_RNO_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \N__3336\,
            in1 => \_gnd_net_\,
            in2 => \N__3310\,
            in3 => \N__3398\,
            lcout => \un1_pulse_len_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_3_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4075\,
            in2 => \_gnd_net_\,
            in3 => \N__3460\,
            lcout => \state_RNIPC4P3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIU5D07_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3399\,
            in2 => \_gnd_net_\,
            in3 => \N__3384\,
            lcout => \state_RNIU5D07\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4103\,
            in2 => \_gnd_net_\,
            in3 => \N__3461\,
            lcout => \state_RNIPC4P3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_8_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3463\,
            in1 => \_gnd_net_\,
            in2 => \N__4115\,
            in3 => \_gnd_net_\,
            lcout => \state_RNIPC4P3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIPC4P3_5_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4104\,
            in2 => \_gnd_net_\,
            in3 => \N__3462\,
            lcout => \state_RNIPC4P3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4822\,
            lcout => \d1.syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI2PCE_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4323\,
            in1 => \N__4338\,
            in2 => \N__4309\,
            in3 => \N__4353\,
            lcout => OPEN,
            ltout => \d1.count_RNI2PCEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI23S21_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3571\,
            in2 => \N__3409\,
            in3 => \_gnd_net_\,
            lcout => \d1.trans_up_1_14\,
            ltout => \d1.trans_up_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI5P873_7_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3535\,
            in1 => \N__3552\,
            in2 => \N__3406\,
            in3 => \N__3541\,
            lcout => s_up,
            ltout => \s_up_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.state_RNIU5D07_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3388\,
            in3 => \N__3383\,
            lcout => \state_RNIU5D07_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI0AFK_16_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3957\,
            in1 => \N__4004\,
            in2 => \N__4522\,
            in3 => \N__4539\,
            lcout => \d1.trans_up_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_RNI5IAP_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__3526\,
            in1 => \N__4554\,
            in2 => \N__3514\,
            in3 => \N__4569\,
            lcout => \d1.trans_up_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNO_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4290\,
            in1 => \N__4251\,
            in2 => \N__4233\,
            in3 => \N__4272\,
            lcout => OPEN,
            ltout => \d1.trans_up_1_13_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_RNO_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3979\,
            in1 => \N__4589\,
            in2 => \N__3565\,
            in3 => \N__4203\,
            lcout => OPEN,
            ltout => \d1.trans_up_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.state_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__3562\,
            in1 => \N__3529\,
            in2 => \N__3556\,
            in3 => \N__3553\,
            lcout => \d1.stateZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNIP9EH_7_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4250\,
            in1 => \N__4271\,
            in2 => \N__4234\,
            in3 => \N__4289\,
            lcout => \d1.trans_up_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_RNI5QJP_11_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4202\,
            in1 => \N__3978\,
            in2 => \N__4591\,
            in3 => \N__3527\,
            lcout => \d1.trans_up_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.sync_1_RNIKI1C_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__3528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3513\,
            lcout => \d1.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3984\,
            in2 => \_gnd_net_\,
            in3 => \N__4008\,
            lcout => \d1.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4794\,
            ce => 'H',
            sr => \N__4506\
        );

    \d1.count_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3983\,
            lcout => \d1.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4794\,
            ce => 'H',
            sr => \N__4506\
        );

    \p.count_RNIL0L01_15_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3938\,
            in1 => \N__3920\,
            in2 => \N__3900\,
            in3 => \N__3875\,
            lcout => \p.count10_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.count_RNIFQK01_12_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3854\,
            in1 => \N__3833\,
            in2 => \N__3814\,
            in3 => \N__3788\,
            lcout => \p.count10_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.count_RNICNK01_10_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3767\,
            in1 => \N__3746\,
            in2 => \N__3727\,
            in3 => \N__3701\,
            lcout => OPEN,
            ltout => \p.count10_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.count_RNIIMK74_10_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3682\,
            in1 => \N__3676\,
            in2 => \N__3670\,
            in3 => \N__3601\,
            lcout => \p.count10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p.count_RNI24M51_1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4459\,
            in1 => \N__3641\,
            in2 => \N__4488\,
            in3 => \N__3620\,
            lcout => \p.count10_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNIE4R8_16_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4870\,
            in1 => \N__4887\,
            in2 => \_gnd_net_\,
            in3 => \N__4731\,
            lcout => \d2.trans_up_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNI6TT21_3_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__4701\,
            in2 => \N__4672\,
            in3 => \N__4716\,
            lcout => \d2.trans_up_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNITE8Q_10_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4623\,
            in1 => \N__4638\,
            in2 => \N__4609\,
            in3 => \N__4653\,
            lcout => \d2.trans_up_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_RNI237_11_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4935\,
            in1 => \N__4950\,
            in2 => \N__4921\,
            in3 => \N__4902\,
            lcout => \d2.count_RNI237Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4159\,
            lcout => \d2.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4138\,
            lcout => \d2.syncZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.sync_1_RNIMV5K_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4129\,
            in2 => \_gnd_net_\,
            in3 => \N__4100\,
            lcout => \d2.idle_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4400\,
            lcout => \d2.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4801\,
            ce => 'H',
            sr => \N__4855\
        );

    \d2.count_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4374\,
            in2 => \_gnd_net_\,
            in3 => \N__4401\,
            lcout => \d2.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4801\,
            ce => 'H',
            sr => \N__4855\
        );

    \d1.un3_count_cry_1_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4009\,
            in2 => \N__3988\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \d1.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d1.count_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3958\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => \d1.countZ0Z_2\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_1\,
            carryout => \d1.un3_count_cry_2\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4354\,
            in2 => \_gnd_net_\,
            in3 => \N__4342\,
            lcout => \d1.countZ0Z_3\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_2\,
            carryout => \d1.un3_count_cry_3\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_4_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4339\,
            in2 => \_gnd_net_\,
            in3 => \N__4327\,
            lcout => \d1.countZ0Z_4\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_3\,
            carryout => \d1.un3_count_cry_4\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_5_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4324\,
            in2 => \_gnd_net_\,
            in3 => \N__4312\,
            lcout => \d1.countZ0Z_5\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_4\,
            carryout => \d1.un3_count_cry_5\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4308\,
            in2 => \_gnd_net_\,
            in3 => \N__4294\,
            lcout => \d1.countZ0Z_6\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_5\,
            carryout => \d1.un3_count_cry_6\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_7_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4291\,
            in2 => \_gnd_net_\,
            in3 => \N__4276\,
            lcout => \d1.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_6\,
            carryout => \d1.un3_count_cry_7\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_8_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4273\,
            in2 => \_gnd_net_\,
            in3 => \N__4255\,
            lcout => \d1.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_7\,
            carryout => \d1.un3_count_cry_8\,
            clk => \N__4799\,
            ce => 'H',
            sr => \N__4507\
        );

    \d1.count_9_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4252\,
            in2 => \_gnd_net_\,
            in3 => \N__4237\,
            lcout => \d1.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \d1.un3_count_cry_9\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_10_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4229\,
            in2 => \_gnd_net_\,
            in3 => \N__4207\,
            lcout => \d1.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_9\,
            carryout => \d1.un3_count_cry_10\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_11_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4204\,
            in2 => \_gnd_net_\,
            in3 => \N__4189\,
            lcout => \d1.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_10\,
            carryout => \d1.un3_count_cry_11\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_12_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4590\,
            in2 => \_gnd_net_\,
            in3 => \N__4573\,
            lcout => \d1.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_11\,
            carryout => \d1.un3_count_cry_12\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_13_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4570\,
            in2 => \_gnd_net_\,
            in3 => \N__4558\,
            lcout => \d1.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_12\,
            carryout => \d1.un3_count_cry_13\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_14_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4555\,
            in2 => \_gnd_net_\,
            in3 => \N__4543\,
            lcout => \d1.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_13\,
            carryout => \d1.un3_count_cry_14\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_15_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4540\,
            in2 => \_gnd_net_\,
            in3 => \N__4528\,
            lcout => \d1.countZ0Z_15\,
            ltout => OPEN,
            carryin => \d1.un3_count_cry_14\,
            carryout => \d1.un3_count_cry_15\,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \d1.count_16_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4521\,
            in2 => \_gnd_net_\,
            in3 => \N__4525\,
            lcout => \d1.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4795\,
            ce => 'H',
            sr => \N__4505\
        );

    \p.count_1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4487\,
            lcout => \p.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4791\,
            ce => \N__4430\,
            sr => \_gnd_net_\
        );

    \p.count_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4463\,
            lcout => \p.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4791\,
            ce => \N__4430\,
            sr => \_gnd_net_\
        );

    \d2.un3_count_cry_1_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4402\,
            in2 => \N__4378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \d2.un3_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d2.count_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4732\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \d2.countZ0Z_2\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_1\,
            carryout => \d2.un3_count_cry_2\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4717\,
            in2 => \_gnd_net_\,
            in3 => \N__4705\,
            lcout => \d2.countZ0Z_3\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_2\,
            carryout => \d2.un3_count_cry_3\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4702\,
            in2 => \_gnd_net_\,
            in3 => \N__4690\,
            lcout => \d2.countZ0Z_4\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_3\,
            carryout => \d2.un3_count_cry_4\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_5_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4687\,
            in2 => \_gnd_net_\,
            in3 => \N__4675\,
            lcout => \d2.countZ0Z_5\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_4\,
            carryout => \d2.un3_count_cry_5\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4671\,
            in2 => \_gnd_net_\,
            in3 => \N__4657\,
            lcout => \d2.countZ0Z_6\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_5\,
            carryout => \d2.un3_count_cry_6\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_7_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4654\,
            in2 => \_gnd_net_\,
            in3 => \N__4642\,
            lcout => \d2.countZ0Z_7\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_6\,
            carryout => \d2.un3_count_cry_7\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_8_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4639\,
            in2 => \_gnd_net_\,
            in3 => \N__4627\,
            lcout => \d2.countZ0Z_8\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_7\,
            carryout => \d2.un3_count_cry_8\,
            clk => \N__4790\,
            ce => 'H',
            sr => \N__4854\
        );

    \d2.count_9_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4624\,
            in2 => \_gnd_net_\,
            in3 => \N__4612\,
            lcout => \d2.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \d2.un3_count_cry_9\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_10_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4605\,
            in2 => \_gnd_net_\,
            in3 => \N__4954\,
            lcout => \d2.countZ0Z_10\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_9\,
            carryout => \d2.un3_count_cry_10\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_11_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4951\,
            in2 => \_gnd_net_\,
            in3 => \N__4939\,
            lcout => \d2.countZ0Z_11\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_10\,
            carryout => \d2.un3_count_cry_11\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_12_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4936\,
            in2 => \_gnd_net_\,
            in3 => \N__4924\,
            lcout => \d2.countZ0Z_12\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_11\,
            carryout => \d2.un3_count_cry_12\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_13_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4920\,
            in2 => \_gnd_net_\,
            in3 => \N__4906\,
            lcout => \d2.countZ0Z_13\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_12\,
            carryout => \d2.un3_count_cry_13\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_14_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4903\,
            in2 => \_gnd_net_\,
            in3 => \N__4891\,
            lcout => \d2.countZ0Z_14\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_13\,
            carryout => \d2.un3_count_cry_14\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_15_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4888\,
            in2 => \_gnd_net_\,
            in3 => \N__4876\,
            lcout => \d2.countZ0Z_15\,
            ltout => OPEN,
            carryin => \d2.un3_count_cry_14\,
            carryout => \d2.un3_count_cry_15\,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d2.count_16_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4869\,
            in2 => \_gnd_net_\,
            in3 => \N__4873\,
            lcout => \d2.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4789\,
            ce => 'H',
            sr => \N__4853\
        );

    \d1.sync_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => \d1.syncZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
