module decoder_7_seg (
  input CLK,
  input [3:0] D,
  output reg [7:0] SEG
  );

always @ ( posedge CLK ) begin

end

endmodule //decoder_7_seg
