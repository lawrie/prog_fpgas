// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Dec 17 2017 21:46:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "timer" view "INTERFACE"

module timer (
    DIGIT,
    SEG2,
    SEG1,
    switch_up,
    switch_start_stop,
    switch_dn,
    switch_cancel,
    CLK,
    BUZZER);

    output [1:0] DIGIT;
    output [7:0] SEG2;
    output [7:0] SEG1;
    input switch_up;
    input switch_start_stop;
    input switch_dn;
    input switch_cancel;
    input CLK;
    output BUZZER;

    wire N__14847;
    wire N__14846;
    wire N__14845;
    wire N__14836;
    wire N__14835;
    wire N__14834;
    wire N__14827;
    wire N__14826;
    wire N__14825;
    wire N__14818;
    wire N__14817;
    wire N__14816;
    wire N__14809;
    wire N__14808;
    wire N__14807;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14791;
    wire N__14790;
    wire N__14789;
    wire N__14782;
    wire N__14781;
    wire N__14780;
    wire N__14773;
    wire N__14772;
    wire N__14771;
    wire N__14764;
    wire N__14763;
    wire N__14762;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14746;
    wire N__14745;
    wire N__14744;
    wire N__14737;
    wire N__14736;
    wire N__14735;
    wire N__14728;
    wire N__14727;
    wire N__14726;
    wire N__14719;
    wire N__14718;
    wire N__14717;
    wire N__14710;
    wire N__14709;
    wire N__14708;
    wire N__14701;
    wire N__14700;
    wire N__14699;
    wire N__14692;
    wire N__14691;
    wire N__14690;
    wire N__14683;
    wire N__14682;
    wire N__14681;
    wire N__14674;
    wire N__14673;
    wire N__14672;
    wire N__14665;
    wire N__14664;
    wire N__14663;
    wire N__14656;
    wire N__14655;
    wire N__14654;
    wire N__14647;
    wire N__14646;
    wire N__14645;
    wire N__14638;
    wire N__14637;
    wire N__14636;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14543;
    wire N__14542;
    wire N__14541;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14524;
    wire N__14523;
    wire N__14522;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14494;
    wire N__14491;
    wire N__14484;
    wire N__14481;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14462;
    wire N__14461;
    wire N__14458;
    wire N__14453;
    wire N__14450;
    wire N__14445;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14424;
    wire N__14423;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14411;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14388;
    wire N__14385;
    wire N__14382;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14360;
    wire N__14357;
    wire N__14352;
    wire N__14351;
    wire N__14350;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14333;
    wire N__14332;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14303;
    wire N__14300;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14276;
    wire N__14275;
    wire N__14274;
    wire N__14273;
    wire N__14272;
    wire N__14271;
    wire N__14270;
    wire N__14269;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14263;
    wire N__14262;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14258;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14250;
    wire N__14249;
    wire N__14248;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14236;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14231;
    wire N__14230;
    wire N__14229;
    wire N__14228;
    wire N__14227;
    wire N__14226;
    wire N__14225;
    wire N__14224;
    wire N__14223;
    wire N__14222;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14216;
    wire N__14215;
    wire N__14214;
    wire N__14213;
    wire N__14212;
    wire N__14211;
    wire N__14210;
    wire N__14209;
    wire N__14208;
    wire N__14207;
    wire N__14206;
    wire N__14205;
    wire N__14204;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14042;
    wire N__14039;
    wire N__14038;
    wire N__14037;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14031;
    wire N__14030;
    wire N__14023;
    wire N__14020;
    wire N__14015;
    wire N__14010;
    wire N__14007;
    wire N__13998;
    wire N__13995;
    wire N__13994;
    wire N__13993;
    wire N__13992;
    wire N__13991;
    wire N__13990;
    wire N__13985;
    wire N__13984;
    wire N__13983;
    wire N__13982;
    wire N__13973;
    wire N__13970;
    wire N__13963;
    wire N__13960;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13868;
    wire N__13867;
    wire N__13866;
    wire N__13863;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13851;
    wire N__13850;
    wire N__13849;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13828;
    wire N__13825;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13794;
    wire N__13791;
    wire N__13790;
    wire N__13789;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13781;
    wire N__13780;
    wire N__13777;
    wire N__13776;
    wire N__13773;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13765;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13757;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13736;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13706;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13680;
    wire N__13679;
    wire N__13676;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13651;
    wire N__13650;
    wire N__13647;
    wire N__13646;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13634;
    wire N__13633;
    wire N__13632;
    wire N__13631;
    wire N__13626;
    wire N__13623;
    wire N__13618;
    wire N__13615;
    wire N__13614;
    wire N__13611;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13585;
    wire N__13582;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13554;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13511;
    wire N__13510;
    wire N__13507;
    wire N__13504;
    wire N__13503;
    wire N__13500;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13489;
    wire N__13488;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13465;
    wire N__13458;
    wire N__13453;
    wire N__13450;
    wire N__13445;
    wire N__13442;
    wire N__13435;
    wire N__13416;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13407;
    wire N__13402;
    wire N__13401;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13386;
    wire N__13383;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13346;
    wire N__13345;
    wire N__13344;
    wire N__13343;
    wire N__13340;
    wire N__13335;
    wire N__13330;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13269;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13257;
    wire N__13254;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13239;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13205;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13143;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13131;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13119;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13074;
    wire N__13073;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13061;
    wire N__13058;
    wire N__13057;
    wire N__13054;
    wire N__13049;
    wire N__13046;
    wire N__13041;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13002;
    wire N__13001;
    wire N__12996;
    wire N__12993;
    wire N__12992;
    wire N__12987;
    wire N__12984;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12965;
    wire N__12960;
    wire N__12957;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12945;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12933;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12918;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12789;
    wire N__12786;
    wire N__12785;
    wire N__12784;
    wire N__12781;
    wire N__12778;
    wire N__12775;
    wire N__12774;
    wire N__12771;
    wire N__12770;
    wire N__12763;
    wire N__12760;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12749;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12732;
    wire N__12731;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12716;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12695;
    wire N__12690;
    wire N__12685;
    wire N__12684;
    wire N__12681;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12642;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12610;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12592;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12576;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12568;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12495;
    wire N__12494;
    wire N__12491;
    wire N__12490;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12468;
    wire N__12465;
    wire N__12456;
    wire N__12453;
    wire N__12452;
    wire N__12451;
    wire N__12450;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12429;
    wire N__12426;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12404;
    wire N__12399;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12367;
    wire N__12362;
    wire N__12357;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12341;
    wire N__12338;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12327;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12315;
    wire N__12310;
    wire N__12305;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12278;
    wire N__12273;
    wire N__12272;
    wire N__12271;
    wire N__12268;
    wire N__12263;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12248;
    wire N__12247;
    wire N__12246;
    wire N__12245;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12228;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12197;
    wire N__12194;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12177;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12156;
    wire N__12155;
    wire N__12152;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12135;
    wire N__12134;
    wire N__12131;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12114;
    wire N__12113;
    wire N__12110;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12100;
    wire N__12097;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12071;
    wire N__12068;
    wire N__12063;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12018;
    wire N__12017;
    wire N__12014;
    wire N__12009;
    wire N__12006;
    wire N__12001;
    wire N__11994;
    wire N__11985;
    wire N__11982;
    wire N__11981;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11969;
    wire N__11964;
    wire N__11959;
    wire N__11958;
    wire N__11955;
    wire N__11950;
    wire N__11949;
    wire N__11946;
    wire N__11945;
    wire N__11940;
    wire N__11933;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11907;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11891;
    wire N__11890;
    wire N__11889;
    wire N__11888;
    wire N__11887;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11878;
    wire N__11873;
    wire N__11870;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11861;
    wire N__11860;
    wire N__11853;
    wire N__11846;
    wire N__11843;
    wire N__11838;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11818;
    wire N__11815;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11794;
    wire N__11791;
    wire N__11784;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11765;
    wire N__11762;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11754;
    wire N__11753;
    wire N__11752;
    wire N__11751;
    wire N__11748;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11728;
    wire N__11725;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11681;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11666;
    wire N__11661;
    wire N__11656;
    wire N__11643;
    wire N__11640;
    wire N__11639;
    wire N__11638;
    wire N__11635;
    wire N__11634;
    wire N__11629;
    wire N__11628;
    wire N__11627;
    wire N__11626;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11609;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11594;
    wire N__11591;
    wire N__11586;
    wire N__11583;
    wire N__11568;
    wire N__11565;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11492;
    wire N__11489;
    wire N__11488;
    wire N__11485;
    wire N__11484;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11459;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11438;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11401;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11299;
    wire N__11294;
    wire N__11291;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11281;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11270;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11238;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11230;
    wire N__11229;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11221;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11181;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11061;
    wire N__11058;
    wire N__11057;
    wire N__11054;
    wire N__11053;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11041;
    wire N__11034;
    wire N__11031;
    wire N__11030;
    wire N__11027;
    wire N__11026;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11014;
    wire N__11007;
    wire N__11006;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10984;
    wire N__10979;
    wire N__10974;
    wire N__10973;
    wire N__10970;
    wire N__10969;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10957;
    wire N__10950;
    wire N__10947;
    wire N__10946;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10919;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10901;
    wire N__10898;
    wire N__10897;
    wire N__10896;
    wire N__10893;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10861;
    wire N__10858;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10826;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10589;
    wire N__10586;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10478;
    wire N__10475;
    wire N__10474;
    wire N__10473;
    wire N__10470;
    wire N__10469;
    wire N__10466;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10446;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10356;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10332;
    wire N__10323;
    wire N__10320;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10289;
    wire N__10288;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10167;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10154;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10136;
    wire N__10125;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10048;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9977;
    wire N__9976;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9941;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9935;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9916;
    wire N__9915;
    wire N__9912;
    wire N__9911;
    wire N__9908;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9870;
    wire N__9869;
    wire N__9868;
    wire N__9867;
    wire N__9866;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9837;
    wire N__9836;
    wire N__9833;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9816;
    wire N__9813;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9789;
    wire N__9786;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9759;
    wire N__9756;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9741;
    wire N__9738;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9657;
    wire N__9654;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9600;
    wire N__9593;
    wire N__9588;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9580;
    wire N__9577;
    wire N__9572;
    wire N__9567;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9555;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9540;
    wire N__9537;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9525;
    wire N__9522;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9486;
    wire N__9483;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9471;
    wire N__9468;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9456;
    wire N__9453;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9441;
    wire N__9438;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9423;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9408;
    wire N__9405;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9390;
    wire N__9387;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9357;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9315;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9303;
    wire N__9300;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9288;
    wire N__9285;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9273;
    wire N__9270;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9153;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9066;
    wire N__9065;
    wire N__9060;
    wire N__9057;
    wire N__9056;
    wire N__9053;
    wire N__9052;
    wire N__9049;
    wire N__9048;
    wire N__9043;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8960;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8934;
    wire N__8933;
    wire N__8930;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8907;
    wire N__8904;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8877;
    wire N__8876;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8850;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8763;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8751;
    wire N__8748;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8635;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8612;
    wire N__8611;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8481;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8469;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8454;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8412;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8400;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8385;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8315;
    wire N__8310;
    wire N__8309;
    wire N__8308;
    wire N__8305;
    wire N__8304;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8289;
    wire N__8280;
    wire N__8277;
    wire N__8276;
    wire N__8271;
    wire N__8270;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8116;
    wire N__8111;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8083;
    wire N__8080;
    wire N__8075;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8057;
    wire N__8056;
    wire N__8055;
    wire N__8054;
    wire N__8053;
    wire N__8052;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8027;
    wire N__8024;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8007;
    wire N__8004;
    wire N__8003;
    wire N__8000;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7983;
    wire N__7980;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7958;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7946;
    wire N__7945;
    wire N__7942;
    wire N__7937;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7891;
    wire N__7886;
    wire N__7883;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7859;
    wire N__7858;
    wire N__7855;
    wire N__7850;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7829;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7784;
    wire N__7783;
    wire N__7780;
    wire N__7775;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7676;
    wire N__7675;
    wire N__7674;
    wire N__7671;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7653;
    wire N__7652;
    wire N__7649;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7632;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7617;
    wire N__7614;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7599;
    wire N__7596;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7584;
    wire N__7581;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7566;
    wire N__7563;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7551;
    wire N__7548;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7509;
    wire N__7506;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7494;
    wire N__7491;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7458;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7431;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7416;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7323;
    wire N__7320;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7308;
    wire N__7305;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7269;
    wire N__7266;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7254;
    wire N__7251;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7239;
    wire N__7236;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7116;
    wire N__7113;
    wire N__7112;
    wire N__7111;
    wire N__7108;
    wire N__7103;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7091;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7079;
    wire N__7074;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7040;
    wire N__7037;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7027;
    wire N__7020;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7008;
    wire N__7005;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6917;
    wire N__6914;
    wire N__6913;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6901;
    wire N__6894;
    wire N__6893;
    wire N__6890;
    wire N__6889;
    wire N__6886;
    wire N__6881;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6866;
    wire N__6865;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6849;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6810;
    wire N__6805;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6771;
    wire N__6758;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6726;
    wire N__6723;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6681;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6669;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6657;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6642;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6528;
    wire N__6525;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6483;
    wire N__6480;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6465;
    wire N__6462;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6447;
    wire N__6444;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6311;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6307;
    wire N__6306;
    wire N__6305;
    wire N__6298;
    wire N__6291;
    wire N__6286;
    wire N__6279;
    wire N__6278;
    wire N__6277;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6256;
    wire N__6255;
    wire N__6254;
    wire N__6249;
    wire N__6246;
    wire N__6241;
    wire N__6234;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6215;
    wire N__6212;
    wire N__6205;
    wire N__6204;
    wire N__6203;
    wire N__6198;
    wire N__6195;
    wire N__6190;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6163;
    wire N__6158;
    wire N__6153;
    wire N__6150;
    wire N__6149;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6126;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6114;
    wire N__6111;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5977;
    wire N__5968;
    wire N__5965;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5936;
    wire N__5935;
    wire N__5932;
    wire N__5931;
    wire N__5930;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5922;
    wire N__5913;
    wire N__5906;
    wire N__5901;
    wire N__5900;
    wire N__5899;
    wire N__5898;
    wire N__5897;
    wire N__5896;
    wire N__5895;
    wire N__5886;
    wire N__5879;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5854;
    wire N__5851;
    wire N__5844;
    wire N__5843;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5829;
    wire N__5822;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire VCCG0;
    wire GNDG0;
    wire SEG1_c_5;
    wire SEG1_c_6;
    wire SEG1_c_4;
    wire SEG1_c_3;
    wire SEG1_c_1;
    wire SEG1_c_2;
    wire SEG1_c_0;
    wire \display1.prescaler8_cascade_ ;
    wire \display1.digit_dataZ0Z_3 ;
    wire DIGIT_c_0;
    wire \display1.digit_dataZ0Z_2 ;
    wire \display1.digit_dataZ0Z_1 ;
    wire \display1.digit_posnZ0 ;
    wire \display1.digit_dataZ0Z_0 ;
    wire \display1.prescaler8 ;
    wire \display1.prescaler8_14 ;
    wire \display1.prescaler8_15_cascade_ ;
    wire \display1.prescaler8_21_cascade_ ;
    wire \display1.prescaler8_17_cascade_ ;
    wire \display1.prescaler8_21 ;
    wire \display1.prescaler8_17 ;
    wire \display1.prescaler8_16 ;
    wire \display1.prescaler8_13 ;
    wire \display1.prescalerZ0Z_1 ;
    wire \display1.prescalerZ0Z_0 ;
    wire bfn_5_13_0_;
    wire \display1.prescalerZ0Z_2 ;
    wire \display1.prescaler_2_cry_1 ;
    wire \display1.prescalerZ0Z_3 ;
    wire \display1.prescaler_2_cry_2 ;
    wire \display1.prescalerZ0Z_4 ;
    wire \display1.prescaler_2_4 ;
    wire \display1.prescaler_2_cry_3 ;
    wire \display1.prescalerZ0Z_5 ;
    wire \display1.prescaler_2_cry_4 ;
    wire \display1.prescalerZ0Z_6 ;
    wire \display1.prescaler_2_6 ;
    wire \display1.prescaler_2_cry_5 ;
    wire \display1.prescalerZ0Z_7 ;
    wire \display1.prescaler_2_cry_6 ;
    wire \display1.prescalerZ0Z_8 ;
    wire \display1.prescaler_2_8 ;
    wire \display1.prescaler_2_cry_7 ;
    wire \display1.prescaler_2_cry_8 ;
    wire \display1.prescalerZ0Z_9 ;
    wire \display1.prescaler_2_9 ;
    wire bfn_5_14_0_;
    wire \display1.prescaler_2_cry_9 ;
    wire \display1.prescaler_2_cry_10 ;
    wire \display1.prescaler_2_cry_11 ;
    wire \display1.prescaler_2_cry_12 ;
    wire \display1.prescalerZ0Z_14 ;
    wire \display1.prescaler_2_14 ;
    wire \display1.prescaler_2_cry_13 ;
    wire \display1.prescalerZ0Z_15 ;
    wire \display1.prescaler_2_15 ;
    wire \display1.prescaler_2_cry_14 ;
    wire \display1.prescalerZ0Z_16 ;
    wire \display1.prescaler_2_cry_15 ;
    wire \display1.prescaler_2_cry_16 ;
    wire \display1.prescalerZ0Z_17 ;
    wire bfn_5_15_0_;
    wire \display1.prescalerZ0Z_18 ;
    wire \display1.prescaler_2_cry_17 ;
    wire \display1.prescalerZ0Z_19 ;
    wire \display1.prescaler_2_cry_18 ;
    wire \display1.prescalerZ0Z_20 ;
    wire \display1.prescaler_2_cry_19 ;
    wire \display1.prescalerZ0Z_21 ;
    wire \display1.prescaler_2_cry_20 ;
    wire \display1.prescalerZ0Z_22 ;
    wire \display1.prescaler_2_cry_21 ;
    wire \display1.prescaler_2_cry_22 ;
    wire \display1.prescalerZ0Z_23 ;
    wire \display1.prescalerZ0Z_12 ;
    wire \display1.prescalerZ0Z_11 ;
    wire \display1.prescalerZ0Z_13 ;
    wire \display1.prescalerZ0Z_10 ;
    wire \display1.prescaler8_12 ;
    wire \d1.idle_i ;
    wire \d1.trans_up_1_11_cascade_ ;
    wire \a.BUZZER3_14_cascade_ ;
    wire \a.BUZZER3_20_cascade_ ;
    wire BUZZER_c;
    wire \a.BUZZER3_20 ;
    wire \a.BUZZER3_19 ;
    wire \a.BUZZER3_18 ;
    wire \a.BUZZER3_17 ;
    wire \a.BUZZER3_16_cascade_ ;
    wire \a.BUZZER3_24 ;
    wire \d1.syncZ0Z_1 ;
    wire \d1.trans_up_1_12_cascade_ ;
    wire \d1.g1_3 ;
    wire \d1.g1_4_cascade_ ;
    wire \d1.countZ0Z_1 ;
    wire bfn_7_16_0_;
    wire \d1.countZ0Z_2 ;
    wire \d1.un3_count_cry_1 ;
    wire \d1.un3_count_cry_2 ;
    wire \d1.un3_count_cry_3 ;
    wire \d1.un3_count_cry_4 ;
    wire \d1.un3_count_cry_5 ;
    wire \d1.un3_count_cry_6 ;
    wire \d1.un3_count_cry_7 ;
    wire \d1.un3_count_cry_8 ;
    wire bfn_7_17_0_;
    wire \d1.un3_count_cry_9 ;
    wire \d1.un3_count_cry_10 ;
    wire \d1.un3_count_cry_11 ;
    wire \d1.countZ0Z_13 ;
    wire \d1.un3_count_cry_12 ;
    wire \d1.countZ0Z_14 ;
    wire \d1.un3_count_cry_13 ;
    wire \d1.countZ0Z_15 ;
    wire \d1.un3_count_cry_14 ;
    wire \d1.un3_count_cry_15 ;
    wire \d1.countZ0Z_16 ;
    wire \d1.idle_i_g ;
    wire switch_dn_c;
    wire \a.countZ0Z_1 ;
    wire bfn_8_11_0_;
    wire \a.countZ0Z_2 ;
    wire \a.count_1_cry_1 ;
    wire \a.countZ0Z_3 ;
    wire \a.count_1_cry_2 ;
    wire \a.countZ0Z_4 ;
    wire \a.count_1_cry_3 ;
    wire \a.countZ0Z_5 ;
    wire \a.count_1_cry_4 ;
    wire \a.countZ0Z_6 ;
    wire \a.count_1_cry_5 ;
    wire \a.countZ0Z_7 ;
    wire \a.count_1_cry_6 ;
    wire \a.countZ0Z_8 ;
    wire \a.count_1_8 ;
    wire \a.count_1_cry_7 ;
    wire \a.count_1_cry_8 ;
    wire \a.countZ0Z_9 ;
    wire bfn_8_12_0_;
    wire \a.countZ0Z_10 ;
    wire \a.count_1_10 ;
    wire \a.count_1_cry_9 ;
    wire \a.countZ0Z_11 ;
    wire \a.count_1_11 ;
    wire \a.count_1_cry_10 ;
    wire \a.countZ0Z_12 ;
    wire \a.count_1_12 ;
    wire \a.count_1_cry_11 ;
    wire \a.countZ0Z_13 ;
    wire \a.count_1_13 ;
    wire \a.count_1_cry_12 ;
    wire \a.countZ0Z_14 ;
    wire \a.count_1_14 ;
    wire \a.count_1_cry_13 ;
    wire \a.countZ0Z_15 ;
    wire \a.count_1_cry_14 ;
    wire \a.countZ0Z_16 ;
    wire \a.count_1_cry_15 ;
    wire \a.count_1_cry_16 ;
    wire \a.countZ0Z_17 ;
    wire bfn_8_13_0_;
    wire \a.count_1_cry_17 ;
    wire \a.count_1_cry_18 ;
    wire \a.count_1_cry_19 ;
    wire \a.count_1_cry_20 ;
    wire \a.countZ0Z_22 ;
    wire \a.count_1_cry_21 ;
    wire \a.countZ0Z_23 ;
    wire \a.count_1_cry_22 ;
    wire \a.countZ0Z_24 ;
    wire \a.count_1_cry_23 ;
    wire \a.count_1_cry_24 ;
    wire bfn_8_14_0_;
    wire \a.countZ0Z_25 ;
    wire \a.countZ0Z_18 ;
    wire \a.countZ0Z_21 ;
    wire \a.countZ0Z_20 ;
    wire \a.countZ0Z_19 ;
    wire \a.BUZZER3_15 ;
    wire prescalerZ0Z_0;
    wire prescalerZ0Z_1;
    wire bfn_8_15_0_;
    wire prescalerZ0Z_2;
    wire prescaler_1_cry_1;
    wire prescalerZ0Z_3;
    wire prescaler_1_cry_2;
    wire prescalerZ0Z_4;
    wire prescaler_1_cry_3;
    wire prescalerZ0Z_5;
    wire prescaler_1_cry_4;
    wire prescalerZ0Z_6;
    wire prescaler_1_cry_5;
    wire prescalerZ0Z_7;
    wire prescaler_1_cry_6;
    wire prescaler_1_cry_7;
    wire prescaler_1_cry_8;
    wire bfn_8_16_0_;
    wire prescaler_1_cry_9;
    wire prescaler_1_cry_10;
    wire prescaler_1_cry_11;
    wire prescaler_1_cry_12;
    wire prescaler_1_cry_13;
    wire prescaler_1_cry_14;
    wire prescaler_1_cry_15;
    wire prescaler_1_cry_16;
    wire bfn_8_17_0_;
    wire prescaler_1_cry_17;
    wire prescaler_1_cry_18;
    wire prescaler_1_cry_19;
    wire prescaler_1_cry_20;
    wire prescaler_1_cry_21;
    wire prescaler_1_cry_22;
    wire prescaler_1_cry_23;
    wire prescaler_1_cry_24;
    wire bfn_8_18_0_;
    wire prescaler_1_cry_25;
    wire prescaler_1_cry_26;
    wire prescaler_1_cry_7_THRU_CO;
    wire prescalerZ0Z_8;
    wire prescaler_1_cry_22_THRU_CO;
    wire prescalerZ0Z_23;
    wire prescaler_1_cry_23_THRU_CO;
    wire prescalerZ0Z_24;
    wire prescaler_1_cry_25_THRU_CO;
    wire prescalerZ0Z_26;
    wire prescaler_1_cry_19_THRU_CO;
    wire prescaler_1_cry_20_THRU_CO;
    wire prescaler_1_cry_21_THRU_CO;
    wire prescaler_1_cry_12_THRU_CO;
    wire prescalerZ0Z_13;
    wire prescaler_1_cry_13_THRU_CO;
    wire prescalerZ0Z_14;
    wire prescaler_1_cry_14_THRU_CO;
    wire prescalerZ0Z_15;
    wire prescaler_1_cry_15_THRU_CO;
    wire prescalerZ0Z_16;
    wire prescaler_1_cry_17_THRU_CO;
    wire un1_state_3_g;
    wire prescalerZ0Z_20;
    wire prescalerZ0Z_21;
    wire prescalerZ0Z_22;
    wire prescalerZ0Z_18;
    wire decrement_time_0_prescaler10_0_and;
    wire bfn_9_13_0_;
    wire decrement_time_0_prescaler10_1_and;
    wire decrement_time_0_prescaler10_0;
    wire decrement_time_0_prescaler10_2_and;
    wire decrement_time_0_prescaler10_1;
    wire decrement_time_0_prescaler10_3_and;
    wire decrement_time_0_prescaler10_2;
    wire decrement_time_0_prescaler10_4_and;
    wire decrement_time_0_prescaler10_3;
    wire decrement_time_0_prescaler10_4;
    wire decrement_time_0_prescaler10_5;
    wire decrement_time_0_prescaler10;
    wire \d1.mins27_1_cascade_ ;
    wire \d1.g2Z0Z_0_cascade_ ;
    wire \d1.g0_1_a5_0_9 ;
    wire \d1.g0_1_a5_0_8 ;
    wire \d1.g0_0_0_a4_2_0 ;
    wire \d1.gZ0Z2 ;
    wire \d1.countZ0Z_0 ;
    wire \d1.countZ0Z_11 ;
    wire \d1.g2_12_0 ;
    wire \d1.g2Z0Z_12_cascade_ ;
    wire prescalerZ0Z_10;
    wire prescalerZ0Z_11;
    wire prescalerZ0Z_9;
    wire prescalerZ0Z_12;
    wire decrement_time_0_prescaler10_5_and;
    wire prescalerZ0Z_25;
    wire prescalerZ0Z_27;
    wire prescalerZ0Z_17;
    wire prescalerZ0Z_19;
    wire decrement_time_0_prescaler10_6_and;
    wire \d1.g2_7_2_cascade_ ;
    wire \d1.countZ0Z_12 ;
    wire switch_cancel_c;
    wire \d3.syncZ0Z_0 ;
    wire \d1.g2_7_1 ;
    wire \d2.syncZ0Z_0 ;
    wire \d4.idle_i ;
    wire \d1.g2Z0Z_1_cascade_ ;
    wire \d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_ ;
    wire \a.countZ0Z_0 ;
    wire \d3.trans_up_1_15_1 ;
    wire \d3.trans_up_1_15_8 ;
    wire \d4.syncZ0Z_1 ;
    wire \d3.trans_up_1_15_7 ;
    wire \d4.trans_up_1_9 ;
    wire \d4.trans_up_1_12 ;
    wire \d4.trans_up_1_11 ;
    wire \d4.trans_up_1_13_cascade_ ;
    wire \d4.trans_up_1_10 ;
    wire d4_trans_up_1_cascade_;
    wire ten_secs_r_1_1_cascade_;
    wire \d3.trans_up_1_14_2_cascade_ ;
    wire s_cancel_cascade_;
    wire d4_state;
    wire d4_trans_up_1;
    wire secs_0_sqmuxa_cascade_;
    wire un1_state_9_0;
    wire \d1.ten_secs_1_sqmuxa_0 ;
    wire \d1.g2_0Z0Z_4 ;
    wire \d1.g2_0Z0Z_3 ;
    wire ten_secs_1_sqmuxa_cascade_;
    wire \d1.g1_0 ;
    wire \d1.g0_0_0_0_0_cascade_ ;
    wire mins_storedZ0Z_1;
    wire \d1.un1_mins_4_0_1_cascade_ ;
    wire \d1.countZ0Z_9 ;
    wire \d1.countZ0Z_8 ;
    wire \d1.countZ0Z_10 ;
    wire \d1.countZ0Z_7 ;
    wire \d1.trans_up_1_9 ;
    wire \d1.g2Z0Z_11 ;
    wire \d1.un1_mins_1_sqmuxa_0_cascade_ ;
    wire \d1.un1_mins_3_sqmuxa_0_0_cascade_ ;
    wire \d1.N_4 ;
    wire mins_storedZ0Z_2;
    wire \d1.g1_cascade_ ;
    wire \d1.g1_7 ;
    wire \d1.g1_8 ;
    wire \d1.g1_14 ;
    wire \d1.g0_1_a5_0_10 ;
    wire \d1.g0_1_a5_0_15 ;
    wire \d1.trans_up_1_10 ;
    wire \d1.trans_up_1_11 ;
    wire \d1.trans_up_1_13 ;
    wire \d1.trans_up_1_0_cascade_ ;
    wire \d1.g0_2_0_o2_2_cascade_ ;
    wire mins_storedZ0Z_0;
    wire \d1.g0_0_0 ;
    wire \d1.N_19_i_cascade_ ;
    wire \d1.stateZ0Z_0 ;
    wire \d1.g2_8_1 ;
    wire \d2.g0_0_10_cascade_ ;
    wire \d2.g0_0_12 ;
    wire \d2.g0_0_14_cascade_ ;
    wire \d1.g2_8_0 ;
    wire \d2.g0_0_11 ;
    wire \d2.trans_up_1_14_2 ;
    wire \d1.g2Z0Z_7_cascade_ ;
    wire \d1.g0_1_0_a4Z0Z_7_cascade_ ;
    wire \d4.countZ0Z_0 ;
    wire \d4.countZ0Z_1 ;
    wire bfn_11_11_0_;
    wire \d4.countZ0Z_2 ;
    wire \d4.un3_count_cry_1 ;
    wire \d4.countZ0Z_3 ;
    wire \d4.un3_count_cry_2 ;
    wire \d4.countZ0Z_4 ;
    wire \d4.un3_count_cry_3 ;
    wire \d4.countZ0Z_5 ;
    wire \d4.un3_count_cry_4 ;
    wire \d4.countZ0Z_6 ;
    wire \d4.un3_count_cry_5 ;
    wire \d4.countZ0Z_7 ;
    wire \d4.un3_count_cry_6 ;
    wire \d4.countZ0Z_8 ;
    wire \d4.un3_count_cry_7 ;
    wire \d4.un3_count_cry_8 ;
    wire \d4.countZ0Z_9 ;
    wire bfn_11_12_0_;
    wire \d4.countZ0Z_10 ;
    wire \d4.un3_count_cry_9 ;
    wire \d4.countZ0Z_11 ;
    wire \d4.un3_count_cry_10 ;
    wire \d4.countZ0Z_12 ;
    wire \d4.un3_count_cry_11 ;
    wire \d4.countZ0Z_13 ;
    wire \d4.un3_count_cry_12 ;
    wire \d4.countZ0Z_14 ;
    wire \d4.un3_count_cry_13 ;
    wire \d4.countZ0Z_15 ;
    wire \d4.un3_count_cry_14 ;
    wire \d4.un3_count_cry_15 ;
    wire \d4.countZ0Z_16 ;
    wire \d4.idle_i_g ;
    wire \d3.countZ0Z_0 ;
    wire \d3.countZ0Z_1 ;
    wire bfn_11_13_0_;
    wire \d3.countZ0Z_2 ;
    wire \d3.un3_count_cry_1 ;
    wire \d3.countZ0Z_3 ;
    wire \d3.un3_count_cry_2 ;
    wire \d3.countZ0Z_4 ;
    wire \d3.un3_count_cry_3 ;
    wire \d3.countZ0Z_5 ;
    wire \d3.un3_count_cry_4 ;
    wire \d3.countZ0Z_6 ;
    wire \d3.un3_count_cry_5 ;
    wire \d3.countZ0Z_7 ;
    wire \d3.un3_count_cry_6 ;
    wire \d3.countZ0Z_8 ;
    wire \d3.un3_count_cry_7 ;
    wire \d3.un3_count_cry_8 ;
    wire \d3.countZ0Z_9 ;
    wire bfn_11_14_0_;
    wire \d3.countZ0Z_10 ;
    wire \d3.un3_count_cry_9 ;
    wire \d3.countZ0Z_11 ;
    wire \d3.un3_count_cry_10 ;
    wire \d3.countZ0Z_12 ;
    wire \d3.un3_count_cry_11 ;
    wire \d3.un3_count_cry_12 ;
    wire \d3.un3_count_cry_13 ;
    wire \d3.un3_count_cry_14 ;
    wire \d3.un3_count_cry_15 ;
    wire \d3.idle_i_g ;
    wire decrement_time_0_prescaler10_THRU_CO;
    wire un1_state_7_0_cascade_;
    wire un1_alarm_on_0_sqmuxa_0_i_cascade_;
    wire N_120_1;
    wire s_cancel;
    wire \d3.countZ0Z_13 ;
    wire d3_g0_1;
    wire \d1.secs_0_sqmuxa_xZ0Z1 ;
    wire mins_storedZ0Z_3;
    wire \d1.N_5 ;
    wire \d1.un1_mins_1_sqmuxa_0 ;
    wire \d1.g0_0_0_a4_2_1 ;
    wire secs_RNO_0Z0Z_2_cascade_;
    wire secs_0_sqmuxa;
    wire un1_state_7_0;
    wire un1_secs_c3_cascade_;
    wire un1_alarm_on_0_sqmuxa_0_i;
    wire \d1.trans_up_1_0 ;
    wire \d1.g2_i_a5_3 ;
    wire \d1.g0_0_0Z0Z_1_cascade_ ;
    wire \d1.g2Z0Z_10 ;
    wire \d1.g0_2_0_a4Z0Z_2 ;
    wire s_dn;
    wire \d1.g0_2_0_o2_2 ;
    wire \d1.g2_i_a5_0Z0Z_3 ;
    wire \d1.g2_i_a5_0Z0Z_6_cascade_ ;
    wire \d1.g2_i_a5Z0Z_2 ;
    wire bfn_11_18_0_;
    wire \d2.un3_count_cry_1 ;
    wire \d2.un3_count_cry_2 ;
    wire \d2.un3_count_cry_3 ;
    wire \d2.un3_count_cry_4 ;
    wire \d2.un3_count_cry_5 ;
    wire \d2.un3_count_cry_6 ;
    wire \d2.un3_count_cry_7 ;
    wire \d2.un3_count_cry_8 ;
    wire bfn_11_19_0_;
    wire \d2.un3_count_cry_9 ;
    wire \d2.un3_count_cry_10 ;
    wire \d2.un3_count_cry_11 ;
    wire \d2.un3_count_cry_12 ;
    wire \d2.un3_count_cry_13 ;
    wire \d2.un3_count_cry_14 ;
    wire \d2.un3_count_cry_15 ;
    wire \d2.idle_i_g ;
    wire un1_state_0_sqmuxa_1_0_0;
    wire \d1.state_1_sqmuxaZ0 ;
    wire un1_state_0_sqmuxa_1_0;
    wire un1_state_0_sqmuxa_1_0_cascade_;
    wire mins_stored_0_sqmuxa;
    wire \d1.state_0_sqmuxaZ0Z_1 ;
    wire \d1.state_0_sqmuxaZ0Z_2 ;
    wire \d1.state_0_sqmuxaZ0Z_2_cascade_ ;
    wire state_0_sqmuxa;
    wire state_0_sqmuxa_cascade_;
    wire alarm_on_0_sqmuxa;
    wire alarm_onZ0;
    wire \d3.countZ0Z_16 ;
    wire \d3.countZ0Z_15 ;
    wire \d3.countZ0Z_14 ;
    wire \d3.count_RNI4GDSZ0Z_16 ;
    wire ten_secsZ0Z_2;
    wire un1_state_3;
    wire \d1.g0_0Z0Z_2 ;
    wire secsZ0Z_2;
    wire secsZ0Z_1;
    wire secsZ0Z_3;
    wire secsZ0Z_0;
    wire decrement_time_0_secs9;
    wire d2_count_6;
    wire d2_count_5;
    wire \d1.g2_7_0_cascade_ ;
    wire \d1.g2_11_0 ;
    wire \d1.N_3 ;
    wire \d3.trans_up_1_14_2 ;
    wire d3_trans_up_1_15;
    wire \d1.countZ0Z_5 ;
    wire \d1.countZ0Z_4 ;
    wire \d1.countZ0Z_6 ;
    wire \d1.countZ0Z_3 ;
    wire \d1.trans_up_1_12 ;
    wire \d1.g1_9_cascade_ ;
    wire \d1.g1_13 ;
    wire un1_alarm_on_0_sqmuxa_0;
    wire \d1.g2_iZ0Z_0 ;
    wire \d1.N_6 ;
    wire ten_secs_1_sqmuxa;
    wire \d1.mins_2_sqmuxa_1 ;
    wire \d1.mins_16_1Z0Z_3 ;
    wire \d1.g3_0_cascade_ ;
    wire \d1.N_8_0 ;
    wire mins_0_sqmuxa;
    wire \d1.g0_1_a5_0Z0Z_11 ;
    wire \d1.g2_12_1 ;
    wire d2_count_4;
    wire d2_count_0;
    wire \d2.trans_up_1_15 ;
    wire \d2.trans_up_1_15_cascade_ ;
    wire s_dn_0;
    wire \d1.g2Z0Z_8 ;
    wire \d1.mins27_0_0 ;
    wire \d1.g2_i_a5_0Z0Z_7 ;
    wire d2_trans_up_1_15_1;
    wire d2_g0_3_cascade_;
    wire \d1.g2_i_a5_1Z0Z_7 ;
    wire \d2.countZ0Z_8 ;
    wire d2_trans_up_1_15_8;
    wire \d2.countZ0Z_9 ;
    wire d2_count_16;
    wire \d2.countZ0Z_10 ;
    wire \d2.countZ0Z_7 ;
    wire \d2.g0_0_13 ;
    wire d2_count_3;
    wire \d1.g2_8_2 ;
    wire \d2.countZ0Z_12 ;
    wire \d2.countZ0Z_13 ;
    wire \d2.countZ0Z_14 ;
    wire \d2.countZ0Z_11 ;
    wire d2_trans_up_1_15_7;
    wire \d1.g2_i_a5_1Z0Z_6 ;
    wire d2_sync_1;
    wire d2_state;
    wire \d2.idle_i ;
    wire d2_g0_3;
    wire \d1.g0_1_0_a4Z0Z_4_cascade_ ;
    wire stateZ0Z_1;
    wire \d1.g0_1_0_a4Z0Z_8 ;
    wire d2_count_15;
    wire d2_count_2;
    wire d2_count_1;
    wire stateZ0Z_0;
    wire d2_g0_1_cascade_;
    wire \d1.g2_i_a5_1Z0Z_3 ;
    wire \d3.syncZ0Z_1 ;
    wire \d3.stateZ0 ;
    wire \d3.idle_i ;
    wire \d1.g0_1_0Z0Z_0 ;
    wire ten_secsZ0Z_1;
    wire ten_secsZ0Z_0;
    wire BNC1;
    wire bfn_14_12_0_;
    wire \display2.prescaler_2_cry_1 ;
    wire \display2.prescaler_2_cry_2 ;
    wire \display2.prescalerZ0Z_4 ;
    wire \display2.prescaler_2_4 ;
    wire \display2.prescaler_2_cry_3 ;
    wire \display2.prescaler_2_cry_4 ;
    wire \display2.prescalerZ0Z_6 ;
    wire \display2.prescaler_2_6 ;
    wire \display2.prescaler_2_cry_5 ;
    wire \display2.prescaler_2_cry_6 ;
    wire \display2.prescalerZ0Z_8 ;
    wire \display2.prescaler_2_8 ;
    wire \display2.prescaler_2_cry_7 ;
    wire \display2.prescaler_2_cry_8 ;
    wire bfn_14_13_0_;
    wire \display2.prescaler_2_cry_9 ;
    wire \display2.prescaler_2_cry_10 ;
    wire \display2.prescaler_2_cry_11 ;
    wire \display2.prescaler_2_cry_12 ;
    wire \display2.prescaler_2_cry_13 ;
    wire \display2.prescaler_2_cry_14 ;
    wire \display2.prescaler_2_cry_15 ;
    wire \display2.prescaler_2_cry_16 ;
    wire bfn_14_14_0_;
    wire \display2.prescaler_2_cry_17 ;
    wire \display2.prescaler_2_cry_18 ;
    wire \display2.prescaler_2_cry_19 ;
    wire \display2.prescaler_2_cry_20 ;
    wire \display2.prescaler_2_cry_21 ;
    wire \display2.prescaler_2_cry_22 ;
    wire \display2.prescalerZ0Z_23 ;
    wire \display2.prescalerZ0Z_21 ;
    wire \display2.prescalerZ0Z_20 ;
    wire \display2.prescalerZ0Z_22 ;
    wire \display2.prescalerZ0Z_19 ;
    wire \display2.prescalerZ0Z_5 ;
    wire \display2.prescalerZ0Z_3 ;
    wire \display2.prescalerZ0Z_7 ;
    wire \display2.prescalerZ0Z_2 ;
    wire \display2.prescalerZ0Z_12 ;
    wire \display2.prescalerZ0Z_10 ;
    wire \display2.prescalerZ0Z_13 ;
    wire \display2.prescalerZ0Z_11 ;
    wire \display2.prescaler8_15 ;
    wire \display2.prescaler8_12_cascade_ ;
    wire \display2.prescaler8_13 ;
    wire \display2.prescaler8_21_cascade_ ;
    wire \display2.prescalerZ0Z_1 ;
    wire \display2.prescaler8_14 ;
    wire \display2.prescaler_2_9 ;
    wire \display2.prescalerZ0Z_9 ;
    wire \display2.prescaler_2_14 ;
    wire \display2.prescalerZ0Z_14 ;
    wire \display2.prescalerZ0Z_17 ;
    wire \display2.prescalerZ0Z_16 ;
    wire \display2.prescalerZ0Z_18 ;
    wire \display2.prescalerZ0Z_0 ;
    wire \display2.prescaler8_17 ;
    wire \display2.prescaler_2_15 ;
    wire \display2.prescaler8_21 ;
    wire \display2.prescaler8_17_cascade_ ;
    wire \display2.prescaler8_16 ;
    wire \display2.prescalerZ0Z_15 ;
    wire switch_up_c;
    wire \d1.syncZ0Z_0 ;
    wire minsZ0Z_3;
    wire minsZ0Z_2;
    wire minsZ0Z_1;
    wire minsZ0Z_0;
    wire \display2.digit_posnZ0 ;
    wire DIGIT_c_1;
    wire \display2.prescaler8 ;
    wire switch_start_stop_c;
    wire \d4.syncZ0Z_0 ;
    wire SEG2_c_0;
    wire SEG2_c_5;
    wire SEG2_c_2;
    wire SEG2_c_1;
    wire SEG2_c_4;
    wire SEG2_c_3;
    wire \display2.digit_dataZ0Z_2 ;
    wire \display2.digit_dataZ0Z_3 ;
    wire \display2.digit_dataZ0Z_1 ;
    wire \display2.digit_dataZ0Z_0 ;
    wire SEG2_c_6;
    wire CLK_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__14845),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__14847),
            .DIN(N__14846),
            .DOUT(N__14845),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__14847),
            .PADOUT(N__14846),
            .PADIN(N__14845),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD BUZZER_obuf_iopad (
            .OE(N__14836),
            .DIN(N__14835),
            .DOUT(N__14834),
            .PACKAGEPIN(BUZZER));
    defparam BUZZER_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUZZER_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUZZER_obuf_preio (
            .PADOEN(N__14836),
            .PADOUT(N__14835),
            .PADIN(N__14834),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__6747),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DIGIT_obuf_0_iopad (
            .OE(N__14827),
            .DIN(N__14826),
            .DOUT(N__14825),
            .PACKAGEPIN(DIGIT[0]));
    defparam DIGIT_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT_obuf_0_preio (
            .PADOEN(N__14827),
            .PADOUT(N__14826),
            .PADIN(N__14825),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5958),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DIGIT_obuf_1_iopad (
            .OE(N__14818),
            .DIN(N__14817),
            .DOUT(N__14816),
            .PACKAGEPIN(DIGIT[1]));
    defparam DIGIT_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT_obuf_1_preio (
            .PADOEN(N__14818),
            .PADOUT(N__14817),
            .PADIN(N__14816),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13374),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_0_iopad (
            .OE(N__14809),
            .DIN(N__14808),
            .DOUT(N__14807),
            .PACKAGEPIN(SEG1[0]));
    defparam SEG1_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_0_preio (
            .PADOEN(N__14809),
            .PADOUT(N__14808),
            .PADIN(N__14807),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__6027),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_1_iopad (
            .OE(N__14800),
            .DIN(N__14799),
            .DOUT(N__14798),
            .PACKAGEPIN(SEG1[1]));
    defparam SEG1_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_1_preio (
            .PADOEN(N__14800),
            .PADOUT(N__14799),
            .PADIN(N__14798),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5763),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_2_iopad (
            .OE(N__14791),
            .DIN(N__14790),
            .DOUT(N__14789),
            .PACKAGEPIN(SEG1[2]));
    defparam SEG1_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_2_preio (
            .PADOEN(N__14791),
            .PADOUT(N__14790),
            .PADIN(N__14789),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__6039),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_3_iopad (
            .OE(N__14782),
            .DIN(N__14781),
            .DOUT(N__14780),
            .PACKAGEPIN(SEG1[3]));
    defparam SEG1_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_3_preio (
            .PADOEN(N__14782),
            .PADOUT(N__14781),
            .PADIN(N__14780),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5772),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_4_iopad (
            .OE(N__14773),
            .DIN(N__14772),
            .DOUT(N__14771),
            .PACKAGEPIN(SEG1[4]));
    defparam SEG1_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_4_preio (
            .PADOEN(N__14773),
            .PADOUT(N__14772),
            .PADIN(N__14771),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5781),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_5_iopad (
            .OE(N__14764),
            .DIN(N__14763),
            .DOUT(N__14762),
            .PACKAGEPIN(SEG1[5]));
    defparam SEG1_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_5_preio (
            .PADOEN(N__14764),
            .PADOUT(N__14763),
            .PADIN(N__14762),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5811),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_6_iopad (
            .OE(N__14755),
            .DIN(N__14754),
            .DOUT(N__14753),
            .PACKAGEPIN(SEG1[6]));
    defparam SEG1_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_6_preio (
            .PADOEN(N__14755),
            .PADOUT(N__14754),
            .PADIN(N__14753),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5796),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG1_obuf_7_iopad (
            .OE(N__14746),
            .DIN(N__14745),
            .DOUT(N__14744),
            .PACKAGEPIN(SEG1[7]));
    defparam SEG1_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam SEG1_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG1_obuf_7_preio (
            .PADOEN(N__14746),
            .PADOUT(N__14745),
            .PADIN(N__14744),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_0_iopad (
            .OE(N__14737),
            .DIN(N__14736),
            .DOUT(N__14735),
            .PACKAGEPIN(SEG2[0]));
    defparam SEG2_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_0_preio (
            .PADOEN(N__14737),
            .PADOUT(N__14736),
            .PADIN(N__14735),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13299),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_1_iopad (
            .OE(N__14728),
            .DIN(N__14727),
            .DOUT(N__14726),
            .PACKAGEPIN(SEG2[1]));
    defparam SEG2_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_1_preio (
            .PADOEN(N__14728),
            .PADOUT(N__14727),
            .PADIN(N__14726),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14589),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_2_iopad (
            .OE(N__14719),
            .DIN(N__14718),
            .DOUT(N__14717),
            .PACKAGEPIN(SEG2[2]));
    defparam SEG2_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_2_preio (
            .PADOEN(N__14719),
            .PADOUT(N__14718),
            .PADIN(N__14717),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14601),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_3_iopad (
            .OE(N__14710),
            .DIN(N__14709),
            .DOUT(N__14708),
            .PACKAGEPIN(SEG2[3]));
    defparam SEG2_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_3_preio (
            .PADOEN(N__14710),
            .PADOUT(N__14709),
            .PADIN(N__14708),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14559),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_4_iopad (
            .OE(N__14701),
            .DIN(N__14700),
            .DOUT(N__14699),
            .PACKAGEPIN(SEG2[4]));
    defparam SEG2_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_4_preio (
            .PADOEN(N__14701),
            .PADOUT(N__14700),
            .PADIN(N__14699),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14574),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_5_iopad (
            .OE(N__14692),
            .DIN(N__14691),
            .DOUT(N__14690),
            .PACKAGEPIN(SEG2[5]));
    defparam SEG2_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_5_preio (
            .PADOEN(N__14692),
            .PADOUT(N__14691),
            .PADIN(N__14690),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14619),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_6_iopad (
            .OE(N__14683),
            .DIN(N__14682),
            .DOUT(N__14681),
            .PACKAGEPIN(SEG2[6]));
    defparam SEG2_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_6_preio (
            .PADOEN(N__14683),
            .PADOUT(N__14682),
            .PADIN(N__14681),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14295),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD SEG2_obuf_7_iopad (
            .OE(N__14674),
            .DIN(N__14673),
            .DOUT(N__14672),
            .PACKAGEPIN(SEG2[7]));
    defparam SEG2_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam SEG2_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO SEG2_obuf_7_preio (
            .PADOEN(N__14674),
            .PADOUT(N__14673),
            .PADIN(N__14672),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_cancel_ibuf_iopad (
            .OE(N__14665),
            .DIN(N__14664),
            .DOUT(N__14663),
            .PACKAGEPIN(switch_cancel));
    defparam switch_cancel_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_cancel_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_cancel_ibuf_preio (
            .PADOEN(N__14665),
            .PADOUT(N__14664),
            .PADIN(N__14663),
            .CLOCKENABLE(),
            .DIN0(switch_cancel_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_dn_ibuf_iopad (
            .OE(N__14656),
            .DIN(N__14655),
            .DOUT(N__14654),
            .PACKAGEPIN(switch_dn));
    defparam switch_dn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_dn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_dn_ibuf_preio (
            .PADOEN(N__14656),
            .PADOUT(N__14655),
            .PADIN(N__14654),
            .CLOCKENABLE(),
            .DIN0(switch_dn_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_start_stop_ibuf_iopad (
            .OE(N__14647),
            .DIN(N__14646),
            .DOUT(N__14645),
            .PACKAGEPIN(switch_start_stop));
    defparam switch_start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_start_stop_ibuf_preio (
            .PADOEN(N__14647),
            .PADOUT(N__14646),
            .PADIN(N__14645),
            .CLOCKENABLE(),
            .DIN0(switch_start_stop_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD switch_up_ibuf_iopad (
            .OE(N__14638),
            .DIN(N__14637),
            .DOUT(N__14636),
            .PACKAGEPIN(switch_up));
    defparam switch_up_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam switch_up_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO switch_up_ibuf_preio (
            .PADOEN(N__14638),
            .PADOUT(N__14637),
            .PADIN(N__14636),
            .CLOCKENABLE(),
            .DIN0(switch_up_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__3446 (
            .O(N__14619),
            .I(N__14616));
    LocalMux I__3445 (
            .O(N__14616),
            .I(N__14613));
    Span4Mux_s2_h I__3444 (
            .O(N__14613),
            .I(N__14610));
    Span4Mux_v I__3443 (
            .O(N__14610),
            .I(N__14607));
    Span4Mux_v I__3442 (
            .O(N__14607),
            .I(N__14604));
    Odrv4 I__3441 (
            .O(N__14604),
            .I(SEG2_c_5));
    IoInMux I__3440 (
            .O(N__14601),
            .I(N__14598));
    LocalMux I__3439 (
            .O(N__14598),
            .I(N__14595));
    Span4Mux_s3_h I__3438 (
            .O(N__14595),
            .I(N__14592));
    Odrv4 I__3437 (
            .O(N__14592),
            .I(SEG2_c_2));
    IoInMux I__3436 (
            .O(N__14589),
            .I(N__14586));
    LocalMux I__3435 (
            .O(N__14586),
            .I(N__14583));
    IoSpan4Mux I__3434 (
            .O(N__14583),
            .I(N__14580));
    Span4Mux_s3_h I__3433 (
            .O(N__14580),
            .I(N__14577));
    Odrv4 I__3432 (
            .O(N__14577),
            .I(SEG2_c_1));
    IoInMux I__3431 (
            .O(N__14574),
            .I(N__14571));
    LocalMux I__3430 (
            .O(N__14571),
            .I(N__14568));
    IoSpan4Mux I__3429 (
            .O(N__14568),
            .I(N__14565));
    Span4Mux_s2_h I__3428 (
            .O(N__14565),
            .I(N__14562));
    Odrv4 I__3427 (
            .O(N__14562),
            .I(SEG2_c_4));
    IoInMux I__3426 (
            .O(N__14559),
            .I(N__14556));
    LocalMux I__3425 (
            .O(N__14556),
            .I(N__14553));
    IoSpan4Mux I__3424 (
            .O(N__14553),
            .I(N__14550));
    Span4Mux_s3_h I__3423 (
            .O(N__14550),
            .I(N__14547));
    Odrv4 I__3422 (
            .O(N__14547),
            .I(SEG2_c_3));
    InMux I__3421 (
            .O(N__14544),
            .I(N__14534));
    InMux I__3420 (
            .O(N__14543),
            .I(N__14534));
    InMux I__3419 (
            .O(N__14542),
            .I(N__14534));
    InMux I__3418 (
            .O(N__14541),
            .I(N__14531));
    LocalMux I__3417 (
            .O(N__14534),
            .I(N__14528));
    LocalMux I__3416 (
            .O(N__14531),
            .I(N__14525));
    Span4Mux_h I__3415 (
            .O(N__14528),
            .I(N__14518));
    Span4Mux_v I__3414 (
            .O(N__14525),
            .I(N__14515));
    InMux I__3413 (
            .O(N__14524),
            .I(N__14510));
    InMux I__3412 (
            .O(N__14523),
            .I(N__14510));
    InMux I__3411 (
            .O(N__14522),
            .I(N__14507));
    CascadeMux I__3410 (
            .O(N__14521),
            .I(N__14504));
    Span4Mux_h I__3409 (
            .O(N__14518),
            .I(N__14501));
    Sp12to4 I__3408 (
            .O(N__14515),
            .I(N__14494));
    LocalMux I__3407 (
            .O(N__14510),
            .I(N__14494));
    LocalMux I__3406 (
            .O(N__14507),
            .I(N__14494));
    InMux I__3405 (
            .O(N__14504),
            .I(N__14491));
    Odrv4 I__3404 (
            .O(N__14501),
            .I(\display2.digit_dataZ0Z_2 ));
    Odrv12 I__3403 (
            .O(N__14494),
            .I(\display2.digit_dataZ0Z_2 ));
    LocalMux I__3402 (
            .O(N__14491),
            .I(\display2.digit_dataZ0Z_2 ));
    CascadeMux I__3401 (
            .O(N__14484),
            .I(N__14481));
    InMux I__3400 (
            .O(N__14481),
            .I(N__14469));
    InMux I__3399 (
            .O(N__14480),
            .I(N__14469));
    InMux I__3398 (
            .O(N__14479),
            .I(N__14469));
    InMux I__3397 (
            .O(N__14478),
            .I(N__14466));
    CascadeMux I__3396 (
            .O(N__14477),
            .I(N__14462));
    InMux I__3395 (
            .O(N__14476),
            .I(N__14458));
    LocalMux I__3394 (
            .O(N__14469),
            .I(N__14453));
    LocalMux I__3393 (
            .O(N__14466),
            .I(N__14453));
    CascadeMux I__3392 (
            .O(N__14465),
            .I(N__14450));
    InMux I__3391 (
            .O(N__14462),
            .I(N__14445));
    InMux I__3390 (
            .O(N__14461),
            .I(N__14445));
    LocalMux I__3389 (
            .O(N__14458),
            .I(N__14440));
    Span4Mux_v I__3388 (
            .O(N__14453),
            .I(N__14440));
    InMux I__3387 (
            .O(N__14450),
            .I(N__14437));
    LocalMux I__3386 (
            .O(N__14445),
            .I(N__14434));
    Span4Mux_h I__3385 (
            .O(N__14440),
            .I(N__14431));
    LocalMux I__3384 (
            .O(N__14437),
            .I(\display2.digit_dataZ0Z_3 ));
    Odrv12 I__3383 (
            .O(N__14434),
            .I(\display2.digit_dataZ0Z_3 ));
    Odrv4 I__3382 (
            .O(N__14431),
            .I(\display2.digit_dataZ0Z_3 ));
    CascadeMux I__3381 (
            .O(N__14424),
            .I(N__14419));
    CascadeMux I__3380 (
            .O(N__14423),
            .I(N__14416));
    InMux I__3379 (
            .O(N__14422),
            .I(N__14411));
    InMux I__3378 (
            .O(N__14419),
            .I(N__14411));
    InMux I__3377 (
            .O(N__14416),
            .I(N__14408));
    LocalMux I__3376 (
            .O(N__14411),
            .I(N__14402));
    LocalMux I__3375 (
            .O(N__14408),
            .I(N__14399));
    CascadeMux I__3374 (
            .O(N__14407),
            .I(N__14396));
    CascadeMux I__3373 (
            .O(N__14406),
            .I(N__14392));
    CascadeMux I__3372 (
            .O(N__14405),
            .I(N__14389));
    Span4Mux_v I__3371 (
            .O(N__14402),
            .I(N__14385));
    Span4Mux_v I__3370 (
            .O(N__14399),
            .I(N__14382));
    InMux I__3369 (
            .O(N__14396),
            .I(N__14375));
    InMux I__3368 (
            .O(N__14395),
            .I(N__14375));
    InMux I__3367 (
            .O(N__14392),
            .I(N__14375));
    InMux I__3366 (
            .O(N__14389),
            .I(N__14372));
    CascadeMux I__3365 (
            .O(N__14388),
            .I(N__14369));
    Sp12to4 I__3364 (
            .O(N__14385),
            .I(N__14360));
    Sp12to4 I__3363 (
            .O(N__14382),
            .I(N__14360));
    LocalMux I__3362 (
            .O(N__14375),
            .I(N__14360));
    LocalMux I__3361 (
            .O(N__14372),
            .I(N__14360));
    InMux I__3360 (
            .O(N__14369),
            .I(N__14357));
    Odrv12 I__3359 (
            .O(N__14360),
            .I(\display2.digit_dataZ0Z_1 ));
    LocalMux I__3358 (
            .O(N__14357),
            .I(\display2.digit_dataZ0Z_1 ));
    InMux I__3357 (
            .O(N__14352),
            .I(N__14345));
    InMux I__3356 (
            .O(N__14351),
            .I(N__14345));
    InMux I__3355 (
            .O(N__14350),
            .I(N__14342));
    LocalMux I__3354 (
            .O(N__14345),
            .I(N__14339));
    LocalMux I__3353 (
            .O(N__14342),
            .I(N__14336));
    Span4Mux_v I__3352 (
            .O(N__14339),
            .I(N__14328));
    Span4Mux_v I__3351 (
            .O(N__14336),
            .I(N__14325));
    InMux I__3350 (
            .O(N__14335),
            .I(N__14318));
    InMux I__3349 (
            .O(N__14334),
            .I(N__14318));
    InMux I__3348 (
            .O(N__14333),
            .I(N__14318));
    InMux I__3347 (
            .O(N__14332),
            .I(N__14315));
    CascadeMux I__3346 (
            .O(N__14331),
            .I(N__14312));
    Sp12to4 I__3345 (
            .O(N__14328),
            .I(N__14303));
    Sp12to4 I__3344 (
            .O(N__14325),
            .I(N__14303));
    LocalMux I__3343 (
            .O(N__14318),
            .I(N__14303));
    LocalMux I__3342 (
            .O(N__14315),
            .I(N__14303));
    InMux I__3341 (
            .O(N__14312),
            .I(N__14300));
    Odrv12 I__3340 (
            .O(N__14303),
            .I(\display2.digit_dataZ0Z_0 ));
    LocalMux I__3339 (
            .O(N__14300),
            .I(\display2.digit_dataZ0Z_0 ));
    IoInMux I__3338 (
            .O(N__14295),
            .I(N__14292));
    LocalMux I__3337 (
            .O(N__14292),
            .I(N__14289));
    Span4Mux_s3_h I__3336 (
            .O(N__14289),
            .I(N__14286));
    Span4Mux_v I__3335 (
            .O(N__14286),
            .I(N__14283));
    Span4Mux_v I__3334 (
            .O(N__14283),
            .I(N__14280));
    Odrv4 I__3333 (
            .O(N__14280),
            .I(SEG2_c_6));
    ClkMux I__3332 (
            .O(N__14277),
            .I(N__14055));
    ClkMux I__3331 (
            .O(N__14276),
            .I(N__14055));
    ClkMux I__3330 (
            .O(N__14275),
            .I(N__14055));
    ClkMux I__3329 (
            .O(N__14274),
            .I(N__14055));
    ClkMux I__3328 (
            .O(N__14273),
            .I(N__14055));
    ClkMux I__3327 (
            .O(N__14272),
            .I(N__14055));
    ClkMux I__3326 (
            .O(N__14271),
            .I(N__14055));
    ClkMux I__3325 (
            .O(N__14270),
            .I(N__14055));
    ClkMux I__3324 (
            .O(N__14269),
            .I(N__14055));
    ClkMux I__3323 (
            .O(N__14268),
            .I(N__14055));
    ClkMux I__3322 (
            .O(N__14267),
            .I(N__14055));
    ClkMux I__3321 (
            .O(N__14266),
            .I(N__14055));
    ClkMux I__3320 (
            .O(N__14265),
            .I(N__14055));
    ClkMux I__3319 (
            .O(N__14264),
            .I(N__14055));
    ClkMux I__3318 (
            .O(N__14263),
            .I(N__14055));
    ClkMux I__3317 (
            .O(N__14262),
            .I(N__14055));
    ClkMux I__3316 (
            .O(N__14261),
            .I(N__14055));
    ClkMux I__3315 (
            .O(N__14260),
            .I(N__14055));
    ClkMux I__3314 (
            .O(N__14259),
            .I(N__14055));
    ClkMux I__3313 (
            .O(N__14258),
            .I(N__14055));
    ClkMux I__3312 (
            .O(N__14257),
            .I(N__14055));
    ClkMux I__3311 (
            .O(N__14256),
            .I(N__14055));
    ClkMux I__3310 (
            .O(N__14255),
            .I(N__14055));
    ClkMux I__3309 (
            .O(N__14254),
            .I(N__14055));
    ClkMux I__3308 (
            .O(N__14253),
            .I(N__14055));
    ClkMux I__3307 (
            .O(N__14252),
            .I(N__14055));
    ClkMux I__3306 (
            .O(N__14251),
            .I(N__14055));
    ClkMux I__3305 (
            .O(N__14250),
            .I(N__14055));
    ClkMux I__3304 (
            .O(N__14249),
            .I(N__14055));
    ClkMux I__3303 (
            .O(N__14248),
            .I(N__14055));
    ClkMux I__3302 (
            .O(N__14247),
            .I(N__14055));
    ClkMux I__3301 (
            .O(N__14246),
            .I(N__14055));
    ClkMux I__3300 (
            .O(N__14245),
            .I(N__14055));
    ClkMux I__3299 (
            .O(N__14244),
            .I(N__14055));
    ClkMux I__3298 (
            .O(N__14243),
            .I(N__14055));
    ClkMux I__3297 (
            .O(N__14242),
            .I(N__14055));
    ClkMux I__3296 (
            .O(N__14241),
            .I(N__14055));
    ClkMux I__3295 (
            .O(N__14240),
            .I(N__14055));
    ClkMux I__3294 (
            .O(N__14239),
            .I(N__14055));
    ClkMux I__3293 (
            .O(N__14238),
            .I(N__14055));
    ClkMux I__3292 (
            .O(N__14237),
            .I(N__14055));
    ClkMux I__3291 (
            .O(N__14236),
            .I(N__14055));
    ClkMux I__3290 (
            .O(N__14235),
            .I(N__14055));
    ClkMux I__3289 (
            .O(N__14234),
            .I(N__14055));
    ClkMux I__3288 (
            .O(N__14233),
            .I(N__14055));
    ClkMux I__3287 (
            .O(N__14232),
            .I(N__14055));
    ClkMux I__3286 (
            .O(N__14231),
            .I(N__14055));
    ClkMux I__3285 (
            .O(N__14230),
            .I(N__14055));
    ClkMux I__3284 (
            .O(N__14229),
            .I(N__14055));
    ClkMux I__3283 (
            .O(N__14228),
            .I(N__14055));
    ClkMux I__3282 (
            .O(N__14227),
            .I(N__14055));
    ClkMux I__3281 (
            .O(N__14226),
            .I(N__14055));
    ClkMux I__3280 (
            .O(N__14225),
            .I(N__14055));
    ClkMux I__3279 (
            .O(N__14224),
            .I(N__14055));
    ClkMux I__3278 (
            .O(N__14223),
            .I(N__14055));
    ClkMux I__3277 (
            .O(N__14222),
            .I(N__14055));
    ClkMux I__3276 (
            .O(N__14221),
            .I(N__14055));
    ClkMux I__3275 (
            .O(N__14220),
            .I(N__14055));
    ClkMux I__3274 (
            .O(N__14219),
            .I(N__14055));
    ClkMux I__3273 (
            .O(N__14218),
            .I(N__14055));
    ClkMux I__3272 (
            .O(N__14217),
            .I(N__14055));
    ClkMux I__3271 (
            .O(N__14216),
            .I(N__14055));
    ClkMux I__3270 (
            .O(N__14215),
            .I(N__14055));
    ClkMux I__3269 (
            .O(N__14214),
            .I(N__14055));
    ClkMux I__3268 (
            .O(N__14213),
            .I(N__14055));
    ClkMux I__3267 (
            .O(N__14212),
            .I(N__14055));
    ClkMux I__3266 (
            .O(N__14211),
            .I(N__14055));
    ClkMux I__3265 (
            .O(N__14210),
            .I(N__14055));
    ClkMux I__3264 (
            .O(N__14209),
            .I(N__14055));
    ClkMux I__3263 (
            .O(N__14208),
            .I(N__14055));
    ClkMux I__3262 (
            .O(N__14207),
            .I(N__14055));
    ClkMux I__3261 (
            .O(N__14206),
            .I(N__14055));
    ClkMux I__3260 (
            .O(N__14205),
            .I(N__14055));
    ClkMux I__3259 (
            .O(N__14204),
            .I(N__14055));
    GlobalMux I__3258 (
            .O(N__14055),
            .I(N__14052));
    gio2CtrlBuf I__3257 (
            .O(N__14052),
            .I(CLK_c_g));
    InMux I__3256 (
            .O(N__14049),
            .I(N__14046));
    LocalMux I__3255 (
            .O(N__14046),
            .I(\display2.prescaler_2_15 ));
    CascadeMux I__3254 (
            .O(N__14043),
            .I(N__14039));
    CascadeMux I__3253 (
            .O(N__14042),
            .I(N__14033));
    InMux I__3252 (
            .O(N__14039),
            .I(N__14023));
    InMux I__3251 (
            .O(N__14038),
            .I(N__14023));
    InMux I__3250 (
            .O(N__14037),
            .I(N__14023));
    InMux I__3249 (
            .O(N__14036),
            .I(N__14020));
    InMux I__3248 (
            .O(N__14033),
            .I(N__14015));
    InMux I__3247 (
            .O(N__14032),
            .I(N__14015));
    InMux I__3246 (
            .O(N__14031),
            .I(N__14010));
    InMux I__3245 (
            .O(N__14030),
            .I(N__14010));
    LocalMux I__3244 (
            .O(N__14023),
            .I(N__14007));
    LocalMux I__3243 (
            .O(N__14020),
            .I(\display2.prescaler8_21 ));
    LocalMux I__3242 (
            .O(N__14015),
            .I(\display2.prescaler8_21 ));
    LocalMux I__3241 (
            .O(N__14010),
            .I(\display2.prescaler8_21 ));
    Odrv4 I__3240 (
            .O(N__14007),
            .I(\display2.prescaler8_21 ));
    CascadeMux I__3239 (
            .O(N__13998),
            .I(\display2.prescaler8_17_cascade_ ));
    InMux I__3238 (
            .O(N__13995),
            .I(N__13985));
    InMux I__3237 (
            .O(N__13994),
            .I(N__13985));
    InMux I__3236 (
            .O(N__13993),
            .I(N__13973));
    InMux I__3235 (
            .O(N__13992),
            .I(N__13973));
    InMux I__3234 (
            .O(N__13991),
            .I(N__13973));
    InMux I__3233 (
            .O(N__13990),
            .I(N__13973));
    LocalMux I__3232 (
            .O(N__13985),
            .I(N__13970));
    InMux I__3231 (
            .O(N__13984),
            .I(N__13963));
    InMux I__3230 (
            .O(N__13983),
            .I(N__13963));
    InMux I__3229 (
            .O(N__13982),
            .I(N__13963));
    LocalMux I__3228 (
            .O(N__13973),
            .I(N__13960));
    Odrv4 I__3227 (
            .O(N__13970),
            .I(\display2.prescaler8_16 ));
    LocalMux I__3226 (
            .O(N__13963),
            .I(\display2.prescaler8_16 ));
    Odrv4 I__3225 (
            .O(N__13960),
            .I(\display2.prescaler8_16 ));
    CascadeMux I__3224 (
            .O(N__13953),
            .I(N__13949));
    InMux I__3223 (
            .O(N__13952),
            .I(N__13946));
    InMux I__3222 (
            .O(N__13949),
            .I(N__13943));
    LocalMux I__3221 (
            .O(N__13946),
            .I(\display2.prescalerZ0Z_15 ));
    LocalMux I__3220 (
            .O(N__13943),
            .I(\display2.prescalerZ0Z_15 ));
    InMux I__3219 (
            .O(N__13938),
            .I(N__13935));
    LocalMux I__3218 (
            .O(N__13935),
            .I(N__13932));
    Span4Mux_v I__3217 (
            .O(N__13932),
            .I(N__13929));
    Sp12to4 I__3216 (
            .O(N__13929),
            .I(N__13926));
    Span12Mux_h I__3215 (
            .O(N__13926),
            .I(N__13923));
    Span12Mux_v I__3214 (
            .O(N__13923),
            .I(N__13920));
    Odrv12 I__3213 (
            .O(N__13920),
            .I(switch_up_c));
    InMux I__3212 (
            .O(N__13917),
            .I(N__13914));
    LocalMux I__3211 (
            .O(N__13914),
            .I(N__13911));
    Span4Mux_v I__3210 (
            .O(N__13911),
            .I(N__13908));
    Span4Mux_h I__3209 (
            .O(N__13908),
            .I(N__13905));
    Span4Mux_h I__3208 (
            .O(N__13905),
            .I(N__13902));
    Odrv4 I__3207 (
            .O(N__13902),
            .I(\d1.syncZ0Z_0 ));
    InMux I__3206 (
            .O(N__13899),
            .I(N__13893));
    InMux I__3205 (
            .O(N__13898),
            .I(N__13889));
    CascadeMux I__3204 (
            .O(N__13897),
            .I(N__13886));
    InMux I__3203 (
            .O(N__13896),
            .I(N__13882));
    LocalMux I__3202 (
            .O(N__13893),
            .I(N__13879));
    InMux I__3201 (
            .O(N__13892),
            .I(N__13876));
    LocalMux I__3200 (
            .O(N__13889),
            .I(N__13873));
    InMux I__3199 (
            .O(N__13886),
            .I(N__13868));
    InMux I__3198 (
            .O(N__13885),
            .I(N__13868));
    LocalMux I__3197 (
            .O(N__13882),
            .I(N__13863));
    Span4Mux_v I__3196 (
            .O(N__13879),
            .I(N__13859));
    LocalMux I__3195 (
            .O(N__13876),
            .I(N__13856));
    Span4Mux_v I__3194 (
            .O(N__13873),
            .I(N__13851));
    LocalMux I__3193 (
            .O(N__13868),
            .I(N__13851));
    InMux I__3192 (
            .O(N__13867),
            .I(N__13845));
    InMux I__3191 (
            .O(N__13866),
            .I(N__13842));
    Span4Mux_h I__3190 (
            .O(N__13863),
            .I(N__13838));
    InMux I__3189 (
            .O(N__13862),
            .I(N__13835));
    Span4Mux_h I__3188 (
            .O(N__13859),
            .I(N__13828));
    Span4Mux_v I__3187 (
            .O(N__13856),
            .I(N__13828));
    Span4Mux_v I__3186 (
            .O(N__13851),
            .I(N__13828));
    InMux I__3185 (
            .O(N__13850),
            .I(N__13825));
    InMux I__3184 (
            .O(N__13849),
            .I(N__13820));
    InMux I__3183 (
            .O(N__13848),
            .I(N__13820));
    LocalMux I__3182 (
            .O(N__13845),
            .I(N__13817));
    LocalMux I__3181 (
            .O(N__13842),
            .I(N__13814));
    InMux I__3180 (
            .O(N__13841),
            .I(N__13811));
    Odrv4 I__3179 (
            .O(N__13838),
            .I(minsZ0Z_3));
    LocalMux I__3178 (
            .O(N__13835),
            .I(minsZ0Z_3));
    Odrv4 I__3177 (
            .O(N__13828),
            .I(minsZ0Z_3));
    LocalMux I__3176 (
            .O(N__13825),
            .I(minsZ0Z_3));
    LocalMux I__3175 (
            .O(N__13820),
            .I(minsZ0Z_3));
    Odrv4 I__3174 (
            .O(N__13817),
            .I(minsZ0Z_3));
    Odrv4 I__3173 (
            .O(N__13814),
            .I(minsZ0Z_3));
    LocalMux I__3172 (
            .O(N__13811),
            .I(minsZ0Z_3));
    InMux I__3171 (
            .O(N__13794),
            .I(N__13791));
    LocalMux I__3170 (
            .O(N__13791),
            .I(N__13785));
    InMux I__3169 (
            .O(N__13790),
            .I(N__13782));
    InMux I__3168 (
            .O(N__13789),
            .I(N__13777));
    InMux I__3167 (
            .O(N__13788),
            .I(N__13773));
    Span4Mux_v I__3166 (
            .O(N__13785),
            .I(N__13769));
    LocalMux I__3165 (
            .O(N__13782),
            .I(N__13766));
    InMux I__3164 (
            .O(N__13781),
            .I(N__13761));
    InMux I__3163 (
            .O(N__13780),
            .I(N__13758));
    LocalMux I__3162 (
            .O(N__13777),
            .I(N__13752));
    InMux I__3161 (
            .O(N__13776),
            .I(N__13749));
    LocalMux I__3160 (
            .O(N__13773),
            .I(N__13744));
    InMux I__3159 (
            .O(N__13772),
            .I(N__13741));
    Span4Mux_h I__3158 (
            .O(N__13769),
            .I(N__13736));
    Span4Mux_v I__3157 (
            .O(N__13766),
            .I(N__13736));
    InMux I__3156 (
            .O(N__13765),
            .I(N__13731));
    InMux I__3155 (
            .O(N__13764),
            .I(N__13731));
    LocalMux I__3154 (
            .O(N__13761),
            .I(N__13728));
    LocalMux I__3153 (
            .O(N__13758),
            .I(N__13725));
    InMux I__3152 (
            .O(N__13757),
            .I(N__13720));
    InMux I__3151 (
            .O(N__13756),
            .I(N__13720));
    InMux I__3150 (
            .O(N__13755),
            .I(N__13717));
    Span4Mux_h I__3149 (
            .O(N__13752),
            .I(N__13714));
    LocalMux I__3148 (
            .O(N__13749),
            .I(N__13711));
    InMux I__3147 (
            .O(N__13748),
            .I(N__13706));
    InMux I__3146 (
            .O(N__13747),
            .I(N__13706));
    Odrv4 I__3145 (
            .O(N__13744),
            .I(minsZ0Z_2));
    LocalMux I__3144 (
            .O(N__13741),
            .I(minsZ0Z_2));
    Odrv4 I__3143 (
            .O(N__13736),
            .I(minsZ0Z_2));
    LocalMux I__3142 (
            .O(N__13731),
            .I(minsZ0Z_2));
    Odrv12 I__3141 (
            .O(N__13728),
            .I(minsZ0Z_2));
    Odrv12 I__3140 (
            .O(N__13725),
            .I(minsZ0Z_2));
    LocalMux I__3139 (
            .O(N__13720),
            .I(minsZ0Z_2));
    LocalMux I__3138 (
            .O(N__13717),
            .I(minsZ0Z_2));
    Odrv4 I__3137 (
            .O(N__13714),
            .I(minsZ0Z_2));
    Odrv4 I__3136 (
            .O(N__13711),
            .I(minsZ0Z_2));
    LocalMux I__3135 (
            .O(N__13706),
            .I(minsZ0Z_2));
    InMux I__3134 (
            .O(N__13683),
            .I(N__13676));
    CascadeMux I__3133 (
            .O(N__13682),
            .I(N__13672));
    CascadeMux I__3132 (
            .O(N__13681),
            .I(N__13667));
    CascadeMux I__3131 (
            .O(N__13680),
            .I(N__13664));
    CascadeMux I__3130 (
            .O(N__13679),
            .I(N__13661));
    LocalMux I__3129 (
            .O(N__13676),
            .I(N__13658));
    InMux I__3128 (
            .O(N__13675),
            .I(N__13655));
    InMux I__3127 (
            .O(N__13672),
            .I(N__13652));
    InMux I__3126 (
            .O(N__13671),
            .I(N__13647));
    InMux I__3125 (
            .O(N__13670),
            .I(N__13641));
    InMux I__3124 (
            .O(N__13667),
            .I(N__13641));
    InMux I__3123 (
            .O(N__13664),
            .I(N__13638));
    InMux I__3122 (
            .O(N__13661),
            .I(N__13635));
    Span4Mux_h I__3121 (
            .O(N__13658),
            .I(N__13626));
    LocalMux I__3120 (
            .O(N__13655),
            .I(N__13626));
    LocalMux I__3119 (
            .O(N__13652),
            .I(N__13623));
    InMux I__3118 (
            .O(N__13651),
            .I(N__13618));
    InMux I__3117 (
            .O(N__13650),
            .I(N__13618));
    LocalMux I__3116 (
            .O(N__13647),
            .I(N__13615));
    CascadeMux I__3115 (
            .O(N__13646),
            .I(N__13611));
    LocalMux I__3114 (
            .O(N__13641),
            .I(N__13604));
    LocalMux I__3113 (
            .O(N__13638),
            .I(N__13604));
    LocalMux I__3112 (
            .O(N__13635),
            .I(N__13604));
    CascadeMux I__3111 (
            .O(N__13634),
            .I(N__13601));
    InMux I__3110 (
            .O(N__13633),
            .I(N__13598));
    InMux I__3109 (
            .O(N__13632),
            .I(N__13595));
    InMux I__3108 (
            .O(N__13631),
            .I(N__13592));
    Span4Mux_h I__3107 (
            .O(N__13626),
            .I(N__13585));
    Span4Mux_h I__3106 (
            .O(N__13623),
            .I(N__13585));
    LocalMux I__3105 (
            .O(N__13618),
            .I(N__13585));
    Span4Mux_h I__3104 (
            .O(N__13615),
            .I(N__13582));
    InMux I__3103 (
            .O(N__13614),
            .I(N__13577));
    InMux I__3102 (
            .O(N__13611),
            .I(N__13577));
    Span4Mux_v I__3101 (
            .O(N__13604),
            .I(N__13574));
    InMux I__3100 (
            .O(N__13601),
            .I(N__13571));
    LocalMux I__3099 (
            .O(N__13598),
            .I(minsZ0Z_1));
    LocalMux I__3098 (
            .O(N__13595),
            .I(minsZ0Z_1));
    LocalMux I__3097 (
            .O(N__13592),
            .I(minsZ0Z_1));
    Odrv4 I__3096 (
            .O(N__13585),
            .I(minsZ0Z_1));
    Odrv4 I__3095 (
            .O(N__13582),
            .I(minsZ0Z_1));
    LocalMux I__3094 (
            .O(N__13577),
            .I(minsZ0Z_1));
    Odrv4 I__3093 (
            .O(N__13574),
            .I(minsZ0Z_1));
    LocalMux I__3092 (
            .O(N__13571),
            .I(minsZ0Z_1));
    InMux I__3091 (
            .O(N__13554),
            .I(N__13551));
    LocalMux I__3090 (
            .O(N__13551),
            .I(N__13539));
    InMux I__3089 (
            .O(N__13550),
            .I(N__13536));
    InMux I__3088 (
            .O(N__13549),
            .I(N__13532));
    CascadeMux I__3087 (
            .O(N__13548),
            .I(N__13529));
    CascadeMux I__3086 (
            .O(N__13547),
            .I(N__13526));
    CascadeMux I__3085 (
            .O(N__13546),
            .I(N__13523));
    InMux I__3084 (
            .O(N__13545),
            .I(N__13518));
    InMux I__3083 (
            .O(N__13544),
            .I(N__13518));
    InMux I__3082 (
            .O(N__13543),
            .I(N__13515));
    InMux I__3081 (
            .O(N__13542),
            .I(N__13512));
    Span4Mux_v I__3080 (
            .O(N__13539),
            .I(N__13507));
    LocalMux I__3079 (
            .O(N__13536),
            .I(N__13504));
    CascadeMux I__3078 (
            .O(N__13535),
            .I(N__13500));
    LocalMux I__3077 (
            .O(N__13532),
            .I(N__13496));
    InMux I__3076 (
            .O(N__13529),
            .I(N__13493));
    InMux I__3075 (
            .O(N__13526),
            .I(N__13490));
    InMux I__3074 (
            .O(N__13523),
            .I(N__13484));
    LocalMux I__3073 (
            .O(N__13518),
            .I(N__13481));
    LocalMux I__3072 (
            .O(N__13515),
            .I(N__13476));
    LocalMux I__3071 (
            .O(N__13512),
            .I(N__13476));
    InMux I__3070 (
            .O(N__13511),
            .I(N__13473));
    InMux I__3069 (
            .O(N__13510),
            .I(N__13470));
    Span4Mux_h I__3068 (
            .O(N__13507),
            .I(N__13465));
    Span4Mux_v I__3067 (
            .O(N__13504),
            .I(N__13465));
    InMux I__3066 (
            .O(N__13503),
            .I(N__13458));
    InMux I__3065 (
            .O(N__13500),
            .I(N__13458));
    InMux I__3064 (
            .O(N__13499),
            .I(N__13458));
    Span4Mux_v I__3063 (
            .O(N__13496),
            .I(N__13453));
    LocalMux I__3062 (
            .O(N__13493),
            .I(N__13453));
    LocalMux I__3061 (
            .O(N__13490),
            .I(N__13450));
    InMux I__3060 (
            .O(N__13489),
            .I(N__13445));
    InMux I__3059 (
            .O(N__13488),
            .I(N__13445));
    InMux I__3058 (
            .O(N__13487),
            .I(N__13442));
    LocalMux I__3057 (
            .O(N__13484),
            .I(N__13435));
    Span4Mux_h I__3056 (
            .O(N__13481),
            .I(N__13435));
    Span4Mux_h I__3055 (
            .O(N__13476),
            .I(N__13435));
    LocalMux I__3054 (
            .O(N__13473),
            .I(minsZ0Z_0));
    LocalMux I__3053 (
            .O(N__13470),
            .I(minsZ0Z_0));
    Odrv4 I__3052 (
            .O(N__13465),
            .I(minsZ0Z_0));
    LocalMux I__3051 (
            .O(N__13458),
            .I(minsZ0Z_0));
    Odrv4 I__3050 (
            .O(N__13453),
            .I(minsZ0Z_0));
    Odrv12 I__3049 (
            .O(N__13450),
            .I(minsZ0Z_0));
    LocalMux I__3048 (
            .O(N__13445),
            .I(minsZ0Z_0));
    LocalMux I__3047 (
            .O(N__13442),
            .I(minsZ0Z_0));
    Odrv4 I__3046 (
            .O(N__13435),
            .I(minsZ0Z_0));
    InMux I__3045 (
            .O(N__13416),
            .I(N__13413));
    LocalMux I__3044 (
            .O(N__13413),
            .I(N__13407));
    InMux I__3043 (
            .O(N__13412),
            .I(N__13402));
    InMux I__3042 (
            .O(N__13411),
            .I(N__13402));
    CascadeMux I__3041 (
            .O(N__13410),
            .I(N__13397));
    Span4Mux_v I__3040 (
            .O(N__13407),
            .I(N__13394));
    LocalMux I__3039 (
            .O(N__13402),
            .I(N__13391));
    InMux I__3038 (
            .O(N__13401),
            .I(N__13386));
    InMux I__3037 (
            .O(N__13400),
            .I(N__13386));
    InMux I__3036 (
            .O(N__13397),
            .I(N__13383));
    Odrv4 I__3035 (
            .O(N__13394),
            .I(\display2.digit_posnZ0 ));
    Odrv4 I__3034 (
            .O(N__13391),
            .I(\display2.digit_posnZ0 ));
    LocalMux I__3033 (
            .O(N__13386),
            .I(\display2.digit_posnZ0 ));
    LocalMux I__3032 (
            .O(N__13383),
            .I(\display2.digit_posnZ0 ));
    IoInMux I__3031 (
            .O(N__13374),
            .I(N__13371));
    LocalMux I__3030 (
            .O(N__13371),
            .I(N__13368));
    IoSpan4Mux I__3029 (
            .O(N__13368),
            .I(N__13365));
    Span4Mux_s2_h I__3028 (
            .O(N__13365),
            .I(N__13362));
    Sp12to4 I__3027 (
            .O(N__13362),
            .I(N__13359));
    Span12Mux_s11_h I__3026 (
            .O(N__13359),
            .I(N__13356));
    Odrv12 I__3025 (
            .O(N__13356),
            .I(DIGIT_c_1));
    CEMux I__3024 (
            .O(N__13353),
            .I(N__13350));
    LocalMux I__3023 (
            .O(N__13350),
            .I(N__13347));
    Span4Mux_h I__3022 (
            .O(N__13347),
            .I(N__13340));
    InMux I__3021 (
            .O(N__13346),
            .I(N__13335));
    InMux I__3020 (
            .O(N__13345),
            .I(N__13335));
    InMux I__3019 (
            .O(N__13344),
            .I(N__13330));
    InMux I__3018 (
            .O(N__13343),
            .I(N__13330));
    Odrv4 I__3017 (
            .O(N__13340),
            .I(\display2.prescaler8 ));
    LocalMux I__3016 (
            .O(N__13335),
            .I(\display2.prescaler8 ));
    LocalMux I__3015 (
            .O(N__13330),
            .I(\display2.prescaler8 ));
    InMux I__3014 (
            .O(N__13323),
            .I(N__13320));
    LocalMux I__3013 (
            .O(N__13320),
            .I(N__13317));
    Span12Mux_h I__3012 (
            .O(N__13317),
            .I(N__13314));
    Odrv12 I__3011 (
            .O(N__13314),
            .I(switch_start_stop_c));
    InMux I__3010 (
            .O(N__13311),
            .I(N__13308));
    LocalMux I__3009 (
            .O(N__13308),
            .I(N__13305));
    Span12Mux_v I__3008 (
            .O(N__13305),
            .I(N__13302));
    Odrv12 I__3007 (
            .O(N__13302),
            .I(\d4.syncZ0Z_0 ));
    IoInMux I__3006 (
            .O(N__13299),
            .I(N__13296));
    LocalMux I__3005 (
            .O(N__13296),
            .I(N__13293));
    Span4Mux_s2_h I__3004 (
            .O(N__13293),
            .I(N__13290));
    Span4Mux_v I__3003 (
            .O(N__13290),
            .I(N__13287));
    Odrv4 I__3002 (
            .O(N__13287),
            .I(SEG2_c_0));
    InMux I__3001 (
            .O(N__13284),
            .I(N__13280));
    InMux I__3000 (
            .O(N__13283),
            .I(N__13277));
    LocalMux I__2999 (
            .O(N__13280),
            .I(N__13274));
    LocalMux I__2998 (
            .O(N__13277),
            .I(\display2.prescalerZ0Z_12 ));
    Odrv4 I__2997 (
            .O(N__13274),
            .I(\display2.prescalerZ0Z_12 ));
    InMux I__2996 (
            .O(N__13269),
            .I(N__13265));
    InMux I__2995 (
            .O(N__13268),
            .I(N__13262));
    LocalMux I__2994 (
            .O(N__13265),
            .I(\display2.prescalerZ0Z_10 ));
    LocalMux I__2993 (
            .O(N__13262),
            .I(\display2.prescalerZ0Z_10 ));
    CascadeMux I__2992 (
            .O(N__13257),
            .I(N__13254));
    InMux I__2991 (
            .O(N__13254),
            .I(N__13250));
    InMux I__2990 (
            .O(N__13253),
            .I(N__13247));
    LocalMux I__2989 (
            .O(N__13250),
            .I(N__13244));
    LocalMux I__2988 (
            .O(N__13247),
            .I(\display2.prescalerZ0Z_13 ));
    Odrv4 I__2987 (
            .O(N__13244),
            .I(\display2.prescalerZ0Z_13 ));
    InMux I__2986 (
            .O(N__13239),
            .I(N__13235));
    InMux I__2985 (
            .O(N__13238),
            .I(N__13232));
    LocalMux I__2984 (
            .O(N__13235),
            .I(\display2.prescalerZ0Z_11 ));
    LocalMux I__2983 (
            .O(N__13232),
            .I(\display2.prescalerZ0Z_11 ));
    InMux I__2982 (
            .O(N__13227),
            .I(N__13224));
    LocalMux I__2981 (
            .O(N__13224),
            .I(N__13221));
    Odrv4 I__2980 (
            .O(N__13221),
            .I(\display2.prescaler8_15 ));
    CascadeMux I__2979 (
            .O(N__13218),
            .I(\display2.prescaler8_12_cascade_ ));
    InMux I__2978 (
            .O(N__13215),
            .I(N__13212));
    LocalMux I__2977 (
            .O(N__13212),
            .I(\display2.prescaler8_13 ));
    CascadeMux I__2976 (
            .O(N__13209),
            .I(\display2.prescaler8_21_cascade_ ));
    CascadeMux I__2975 (
            .O(N__13206),
            .I(N__13201));
    InMux I__2974 (
            .O(N__13205),
            .I(N__13198));
    InMux I__2973 (
            .O(N__13204),
            .I(N__13195));
    InMux I__2972 (
            .O(N__13201),
            .I(N__13192));
    LocalMux I__2971 (
            .O(N__13198),
            .I(\display2.prescalerZ0Z_1 ));
    LocalMux I__2970 (
            .O(N__13195),
            .I(\display2.prescalerZ0Z_1 ));
    LocalMux I__2969 (
            .O(N__13192),
            .I(\display2.prescalerZ0Z_1 ));
    InMux I__2968 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__2967 (
            .O(N__13182),
            .I(\display2.prescaler8_14 ));
    InMux I__2966 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__2965 (
            .O(N__13176),
            .I(\display2.prescaler_2_9 ));
    InMux I__2964 (
            .O(N__13173),
            .I(N__13169));
    InMux I__2963 (
            .O(N__13172),
            .I(N__13166));
    LocalMux I__2962 (
            .O(N__13169),
            .I(\display2.prescalerZ0Z_9 ));
    LocalMux I__2961 (
            .O(N__13166),
            .I(\display2.prescalerZ0Z_9 ));
    InMux I__2960 (
            .O(N__13161),
            .I(N__13158));
    LocalMux I__2959 (
            .O(N__13158),
            .I(\display2.prescaler_2_14 ));
    InMux I__2958 (
            .O(N__13155),
            .I(N__13151));
    InMux I__2957 (
            .O(N__13154),
            .I(N__13148));
    LocalMux I__2956 (
            .O(N__13151),
            .I(\display2.prescalerZ0Z_14 ));
    LocalMux I__2955 (
            .O(N__13148),
            .I(\display2.prescalerZ0Z_14 ));
    InMux I__2954 (
            .O(N__13143),
            .I(N__13139));
    InMux I__2953 (
            .O(N__13142),
            .I(N__13136));
    LocalMux I__2952 (
            .O(N__13139),
            .I(\display2.prescalerZ0Z_17 ));
    LocalMux I__2951 (
            .O(N__13136),
            .I(\display2.prescalerZ0Z_17 ));
    InMux I__2950 (
            .O(N__13131),
            .I(N__13127));
    InMux I__2949 (
            .O(N__13130),
            .I(N__13124));
    LocalMux I__2948 (
            .O(N__13127),
            .I(\display2.prescalerZ0Z_16 ));
    LocalMux I__2947 (
            .O(N__13124),
            .I(\display2.prescalerZ0Z_16 ));
    CascadeMux I__2946 (
            .O(N__13119),
            .I(N__13115));
    InMux I__2945 (
            .O(N__13118),
            .I(N__13112));
    InMux I__2944 (
            .O(N__13115),
            .I(N__13109));
    LocalMux I__2943 (
            .O(N__13112),
            .I(\display2.prescalerZ0Z_18 ));
    LocalMux I__2942 (
            .O(N__13109),
            .I(\display2.prescalerZ0Z_18 ));
    InMux I__2941 (
            .O(N__13104),
            .I(N__13096));
    InMux I__2940 (
            .O(N__13103),
            .I(N__13096));
    InMux I__2939 (
            .O(N__13102),
            .I(N__13093));
    InMux I__2938 (
            .O(N__13101),
            .I(N__13090));
    LocalMux I__2937 (
            .O(N__13096),
            .I(\display2.prescalerZ0Z_0 ));
    LocalMux I__2936 (
            .O(N__13093),
            .I(\display2.prescalerZ0Z_0 ));
    LocalMux I__2935 (
            .O(N__13090),
            .I(\display2.prescalerZ0Z_0 ));
    CascadeMux I__2934 (
            .O(N__13083),
            .I(N__13078));
    CascadeMux I__2933 (
            .O(N__13082),
            .I(N__13075));
    CascadeMux I__2932 (
            .O(N__13081),
            .I(N__13070));
    InMux I__2931 (
            .O(N__13078),
            .I(N__13061));
    InMux I__2930 (
            .O(N__13075),
            .I(N__13061));
    InMux I__2929 (
            .O(N__13074),
            .I(N__13061));
    CascadeMux I__2928 (
            .O(N__13073),
            .I(N__13058));
    InMux I__2927 (
            .O(N__13070),
            .I(N__13054));
    InMux I__2926 (
            .O(N__13069),
            .I(N__13049));
    InMux I__2925 (
            .O(N__13068),
            .I(N__13049));
    LocalMux I__2924 (
            .O(N__13061),
            .I(N__13046));
    InMux I__2923 (
            .O(N__13058),
            .I(N__13041));
    InMux I__2922 (
            .O(N__13057),
            .I(N__13041));
    LocalMux I__2921 (
            .O(N__13054),
            .I(\display2.prescaler8_17 ));
    LocalMux I__2920 (
            .O(N__13049),
            .I(\display2.prescaler8_17 ));
    Odrv4 I__2919 (
            .O(N__13046),
            .I(\display2.prescaler8_17 ));
    LocalMux I__2918 (
            .O(N__13041),
            .I(\display2.prescaler8_17 ));
    InMux I__2917 (
            .O(N__13032),
            .I(\display2.prescaler_2_cry_18 ));
    InMux I__2916 (
            .O(N__13029),
            .I(\display2.prescaler_2_cry_19 ));
    InMux I__2915 (
            .O(N__13026),
            .I(\display2.prescaler_2_cry_20 ));
    InMux I__2914 (
            .O(N__13023),
            .I(\display2.prescaler_2_cry_21 ));
    InMux I__2913 (
            .O(N__13020),
            .I(\display2.prescaler_2_cry_22 ));
    CascadeMux I__2912 (
            .O(N__13017),
            .I(N__13013));
    InMux I__2911 (
            .O(N__13016),
            .I(N__13010));
    InMux I__2910 (
            .O(N__13013),
            .I(N__13007));
    LocalMux I__2909 (
            .O(N__13010),
            .I(\display2.prescalerZ0Z_23 ));
    LocalMux I__2908 (
            .O(N__13007),
            .I(\display2.prescalerZ0Z_23 ));
    InMux I__2907 (
            .O(N__13002),
            .I(N__12996));
    InMux I__2906 (
            .O(N__13001),
            .I(N__12996));
    LocalMux I__2905 (
            .O(N__12996),
            .I(\display2.prescalerZ0Z_21 ));
    InMux I__2904 (
            .O(N__12993),
            .I(N__12987));
    InMux I__2903 (
            .O(N__12992),
            .I(N__12987));
    LocalMux I__2902 (
            .O(N__12987),
            .I(\display2.prescalerZ0Z_20 ));
    CascadeMux I__2901 (
            .O(N__12984),
            .I(N__12980));
    CascadeMux I__2900 (
            .O(N__12983),
            .I(N__12977));
    InMux I__2899 (
            .O(N__12980),
            .I(N__12972));
    InMux I__2898 (
            .O(N__12977),
            .I(N__12972));
    LocalMux I__2897 (
            .O(N__12972),
            .I(\display2.prescalerZ0Z_22 ));
    CascadeMux I__2896 (
            .O(N__12969),
            .I(N__12966));
    InMux I__2895 (
            .O(N__12966),
            .I(N__12960));
    InMux I__2894 (
            .O(N__12965),
            .I(N__12960));
    LocalMux I__2893 (
            .O(N__12960),
            .I(\display2.prescalerZ0Z_19 ));
    InMux I__2892 (
            .O(N__12957),
            .I(N__12953));
    InMux I__2891 (
            .O(N__12956),
            .I(N__12950));
    LocalMux I__2890 (
            .O(N__12953),
            .I(\display2.prescalerZ0Z_5 ));
    LocalMux I__2889 (
            .O(N__12950),
            .I(\display2.prescalerZ0Z_5 ));
    InMux I__2888 (
            .O(N__12945),
            .I(N__12941));
    InMux I__2887 (
            .O(N__12944),
            .I(N__12938));
    LocalMux I__2886 (
            .O(N__12941),
            .I(\display2.prescalerZ0Z_3 ));
    LocalMux I__2885 (
            .O(N__12938),
            .I(\display2.prescalerZ0Z_3 ));
    CascadeMux I__2884 (
            .O(N__12933),
            .I(N__12929));
    InMux I__2883 (
            .O(N__12932),
            .I(N__12926));
    InMux I__2882 (
            .O(N__12929),
            .I(N__12923));
    LocalMux I__2881 (
            .O(N__12926),
            .I(\display2.prescalerZ0Z_7 ));
    LocalMux I__2880 (
            .O(N__12923),
            .I(\display2.prescalerZ0Z_7 ));
    InMux I__2879 (
            .O(N__12918),
            .I(N__12914));
    InMux I__2878 (
            .O(N__12917),
            .I(N__12911));
    LocalMux I__2877 (
            .O(N__12914),
            .I(\display2.prescalerZ0Z_2 ));
    LocalMux I__2876 (
            .O(N__12911),
            .I(\display2.prescalerZ0Z_2 ));
    InMux I__2875 (
            .O(N__12906),
            .I(\display2.prescaler_2_cry_9 ));
    InMux I__2874 (
            .O(N__12903),
            .I(\display2.prescaler_2_cry_10 ));
    InMux I__2873 (
            .O(N__12900),
            .I(\display2.prescaler_2_cry_11 ));
    InMux I__2872 (
            .O(N__12897),
            .I(\display2.prescaler_2_cry_12 ));
    InMux I__2871 (
            .O(N__12894),
            .I(\display2.prescaler_2_cry_13 ));
    InMux I__2870 (
            .O(N__12891),
            .I(\display2.prescaler_2_cry_14 ));
    InMux I__2869 (
            .O(N__12888),
            .I(\display2.prescaler_2_cry_15 ));
    InMux I__2868 (
            .O(N__12885),
            .I(bfn_14_14_0_));
    InMux I__2867 (
            .O(N__12882),
            .I(\display2.prescaler_2_cry_17 ));
    InMux I__2866 (
            .O(N__12879),
            .I(\display2.prescaler_2_cry_1 ));
    InMux I__2865 (
            .O(N__12876),
            .I(\display2.prescaler_2_cry_2 ));
    InMux I__2864 (
            .O(N__12873),
            .I(N__12869));
    InMux I__2863 (
            .O(N__12872),
            .I(N__12866));
    LocalMux I__2862 (
            .O(N__12869),
            .I(\display2.prescalerZ0Z_4 ));
    LocalMux I__2861 (
            .O(N__12866),
            .I(\display2.prescalerZ0Z_4 ));
    InMux I__2860 (
            .O(N__12861),
            .I(N__12858));
    LocalMux I__2859 (
            .O(N__12858),
            .I(\display2.prescaler_2_4 ));
    InMux I__2858 (
            .O(N__12855),
            .I(\display2.prescaler_2_cry_3 ));
    InMux I__2857 (
            .O(N__12852),
            .I(\display2.prescaler_2_cry_4 ));
    InMux I__2856 (
            .O(N__12849),
            .I(N__12845));
    InMux I__2855 (
            .O(N__12848),
            .I(N__12842));
    LocalMux I__2854 (
            .O(N__12845),
            .I(\display2.prescalerZ0Z_6 ));
    LocalMux I__2853 (
            .O(N__12842),
            .I(\display2.prescalerZ0Z_6 ));
    InMux I__2852 (
            .O(N__12837),
            .I(N__12834));
    LocalMux I__2851 (
            .O(N__12834),
            .I(\display2.prescaler_2_6 ));
    InMux I__2850 (
            .O(N__12831),
            .I(\display2.prescaler_2_cry_5 ));
    InMux I__2849 (
            .O(N__12828),
            .I(\display2.prescaler_2_cry_6 ));
    InMux I__2848 (
            .O(N__12825),
            .I(N__12821));
    InMux I__2847 (
            .O(N__12824),
            .I(N__12818));
    LocalMux I__2846 (
            .O(N__12821),
            .I(\display2.prescalerZ0Z_8 ));
    LocalMux I__2845 (
            .O(N__12818),
            .I(\display2.prescalerZ0Z_8 ));
    InMux I__2844 (
            .O(N__12813),
            .I(N__12810));
    LocalMux I__2843 (
            .O(N__12810),
            .I(\display2.prescaler_2_8 ));
    InMux I__2842 (
            .O(N__12807),
            .I(\display2.prescaler_2_cry_7 ));
    InMux I__2841 (
            .O(N__12804),
            .I(bfn_14_13_0_));
    CascadeMux I__2840 (
            .O(N__12801),
            .I(N__12792));
    CascadeMux I__2839 (
            .O(N__12800),
            .I(N__12786));
    CascadeMux I__2838 (
            .O(N__12799),
            .I(N__12781));
    InMux I__2837 (
            .O(N__12798),
            .I(N__12778));
    CascadeMux I__2836 (
            .O(N__12797),
            .I(N__12775));
    CascadeMux I__2835 (
            .O(N__12796),
            .I(N__12771));
    InMux I__2834 (
            .O(N__12795),
            .I(N__12763));
    InMux I__2833 (
            .O(N__12792),
            .I(N__12763));
    InMux I__2832 (
            .O(N__12791),
            .I(N__12763));
    InMux I__2831 (
            .O(N__12790),
            .I(N__12760));
    InMux I__2830 (
            .O(N__12789),
            .I(N__12756));
    InMux I__2829 (
            .O(N__12786),
            .I(N__12753));
    InMux I__2828 (
            .O(N__12785),
            .I(N__12750));
    InMux I__2827 (
            .O(N__12784),
            .I(N__12745));
    InMux I__2826 (
            .O(N__12781),
            .I(N__12742));
    LocalMux I__2825 (
            .O(N__12778),
            .I(N__12739));
    InMux I__2824 (
            .O(N__12775),
            .I(N__12736));
    InMux I__2823 (
            .O(N__12774),
            .I(N__12733));
    InMux I__2822 (
            .O(N__12771),
            .I(N__12726));
    InMux I__2821 (
            .O(N__12770),
            .I(N__12726));
    LocalMux I__2820 (
            .O(N__12763),
            .I(N__12723));
    LocalMux I__2819 (
            .O(N__12760),
            .I(N__12720));
    InMux I__2818 (
            .O(N__12759),
            .I(N__12717));
    LocalMux I__2817 (
            .O(N__12756),
            .I(N__12709));
    LocalMux I__2816 (
            .O(N__12753),
            .I(N__12709));
    LocalMux I__2815 (
            .O(N__12750),
            .I(N__12709));
    InMux I__2814 (
            .O(N__12749),
            .I(N__12706));
    InMux I__2813 (
            .O(N__12748),
            .I(N__12703));
    LocalMux I__2812 (
            .O(N__12745),
            .I(N__12700));
    LocalMux I__2811 (
            .O(N__12742),
            .I(N__12695));
    Span4Mux_h I__2810 (
            .O(N__12739),
            .I(N__12695));
    LocalMux I__2809 (
            .O(N__12736),
            .I(N__12690));
    LocalMux I__2808 (
            .O(N__12733),
            .I(N__12690));
    InMux I__2807 (
            .O(N__12732),
            .I(N__12685));
    InMux I__2806 (
            .O(N__12731),
            .I(N__12685));
    LocalMux I__2805 (
            .O(N__12726),
            .I(N__12681));
    Span4Mux_h I__2804 (
            .O(N__12723),
            .I(N__12676));
    Span4Mux_h I__2803 (
            .O(N__12720),
            .I(N__12676));
    LocalMux I__2802 (
            .O(N__12717),
            .I(N__12673));
    InMux I__2801 (
            .O(N__12716),
            .I(N__12670));
    Span4Mux_v I__2800 (
            .O(N__12709),
            .I(N__12667));
    LocalMux I__2799 (
            .O(N__12706),
            .I(N__12656));
    LocalMux I__2798 (
            .O(N__12703),
            .I(N__12656));
    Span4Mux_v I__2797 (
            .O(N__12700),
            .I(N__12656));
    Span4Mux_h I__2796 (
            .O(N__12695),
            .I(N__12656));
    Span4Mux_v I__2795 (
            .O(N__12690),
            .I(N__12656));
    LocalMux I__2794 (
            .O(N__12685),
            .I(N__12653));
    InMux I__2793 (
            .O(N__12684),
            .I(N__12650));
    Span4Mux_h I__2792 (
            .O(N__12681),
            .I(N__12647));
    Span4Mux_v I__2791 (
            .O(N__12676),
            .I(N__12642));
    Span4Mux_h I__2790 (
            .O(N__12673),
            .I(N__12642));
    LocalMux I__2789 (
            .O(N__12670),
            .I(stateZ0Z_0));
    Odrv4 I__2788 (
            .O(N__12667),
            .I(stateZ0Z_0));
    Odrv4 I__2787 (
            .O(N__12656),
            .I(stateZ0Z_0));
    Odrv12 I__2786 (
            .O(N__12653),
            .I(stateZ0Z_0));
    LocalMux I__2785 (
            .O(N__12650),
            .I(stateZ0Z_0));
    Odrv4 I__2784 (
            .O(N__12647),
            .I(stateZ0Z_0));
    Odrv4 I__2783 (
            .O(N__12642),
            .I(stateZ0Z_0));
    CascadeMux I__2782 (
            .O(N__12627),
            .I(d2_g0_1_cascade_));
    InMux I__2781 (
            .O(N__12624),
            .I(N__12621));
    LocalMux I__2780 (
            .O(N__12621),
            .I(\d1.g2_i_a5_1Z0Z_3 ));
    InMux I__2779 (
            .O(N__12618),
            .I(N__12614));
    CascadeMux I__2778 (
            .O(N__12617),
            .I(N__12611));
    LocalMux I__2777 (
            .O(N__12614),
            .I(N__12606));
    InMux I__2776 (
            .O(N__12611),
            .I(N__12603));
    InMux I__2775 (
            .O(N__12610),
            .I(N__12600));
    InMux I__2774 (
            .O(N__12609),
            .I(N__12597));
    Span4Mux_v I__2773 (
            .O(N__12606),
            .I(N__12592));
    LocalMux I__2772 (
            .O(N__12603),
            .I(N__12592));
    LocalMux I__2771 (
            .O(N__12600),
            .I(N__12587));
    LocalMux I__2770 (
            .O(N__12597),
            .I(N__12587));
    Span4Mux_h I__2769 (
            .O(N__12592),
            .I(N__12584));
    Span4Mux_h I__2768 (
            .O(N__12587),
            .I(N__12581));
    Odrv4 I__2767 (
            .O(N__12584),
            .I(\d3.syncZ0Z_1 ));
    Odrv4 I__2766 (
            .O(N__12581),
            .I(\d3.syncZ0Z_1 ));
    InMux I__2765 (
            .O(N__12576),
            .I(N__12572));
    InMux I__2764 (
            .O(N__12575),
            .I(N__12569));
    LocalMux I__2763 (
            .O(N__12572),
            .I(N__12564));
    LocalMux I__2762 (
            .O(N__12569),
            .I(N__12561));
    InMux I__2761 (
            .O(N__12568),
            .I(N__12558));
    InMux I__2760 (
            .O(N__12567),
            .I(N__12555));
    Span4Mux_h I__2759 (
            .O(N__12564),
            .I(N__12552));
    Odrv4 I__2758 (
            .O(N__12561),
            .I(\d3.stateZ0 ));
    LocalMux I__2757 (
            .O(N__12558),
            .I(\d3.stateZ0 ));
    LocalMux I__2756 (
            .O(N__12555),
            .I(\d3.stateZ0 ));
    Odrv4 I__2755 (
            .O(N__12552),
            .I(\d3.stateZ0 ));
    IoInMux I__2754 (
            .O(N__12543),
            .I(N__12540));
    LocalMux I__2753 (
            .O(N__12540),
            .I(N__12537));
    Span4Mux_s2_h I__2752 (
            .O(N__12537),
            .I(N__12534));
    Span4Mux_h I__2751 (
            .O(N__12534),
            .I(N__12531));
    Span4Mux_h I__2750 (
            .O(N__12531),
            .I(N__12528));
    Span4Mux_h I__2749 (
            .O(N__12528),
            .I(N__12525));
    Odrv4 I__2748 (
            .O(N__12525),
            .I(\d3.idle_i ));
    CascadeMux I__2747 (
            .O(N__12522),
            .I(N__12519));
    InMux I__2746 (
            .O(N__12519),
            .I(N__12516));
    LocalMux I__2745 (
            .O(N__12516),
            .I(N__12513));
    Span4Mux_v I__2744 (
            .O(N__12513),
            .I(N__12510));
    Odrv4 I__2743 (
            .O(N__12510),
            .I(\d1.g0_1_0Z0Z_0 ));
    InMux I__2742 (
            .O(N__12507),
            .I(N__12502));
    InMux I__2741 (
            .O(N__12506),
            .I(N__12499));
    InMux I__2740 (
            .O(N__12505),
            .I(N__12496));
    LocalMux I__2739 (
            .O(N__12502),
            .I(N__12491));
    LocalMux I__2738 (
            .O(N__12499),
            .I(N__12485));
    LocalMux I__2737 (
            .O(N__12496),
            .I(N__12485));
    InMux I__2736 (
            .O(N__12495),
            .I(N__12482));
    InMux I__2735 (
            .O(N__12494),
            .I(N__12479));
    Span12Mux_h I__2734 (
            .O(N__12491),
            .I(N__12476));
    InMux I__2733 (
            .O(N__12490),
            .I(N__12473));
    Span4Mux_v I__2732 (
            .O(N__12485),
            .I(N__12468));
    LocalMux I__2731 (
            .O(N__12482),
            .I(N__12468));
    LocalMux I__2730 (
            .O(N__12479),
            .I(N__12465));
    Odrv12 I__2729 (
            .O(N__12476),
            .I(ten_secsZ0Z_1));
    LocalMux I__2728 (
            .O(N__12473),
            .I(ten_secsZ0Z_1));
    Odrv4 I__2727 (
            .O(N__12468),
            .I(ten_secsZ0Z_1));
    Odrv4 I__2726 (
            .O(N__12465),
            .I(ten_secsZ0Z_1));
    InMux I__2725 (
            .O(N__12456),
            .I(N__12453));
    LocalMux I__2724 (
            .O(N__12453),
            .I(N__12446));
    InMux I__2723 (
            .O(N__12452),
            .I(N__12443));
    InMux I__2722 (
            .O(N__12451),
            .I(N__12440));
    InMux I__2721 (
            .O(N__12450),
            .I(N__12437));
    InMux I__2720 (
            .O(N__12449),
            .I(N__12433));
    Span4Mux_h I__2719 (
            .O(N__12446),
            .I(N__12430));
    LocalMux I__2718 (
            .O(N__12443),
            .I(N__12426));
    LocalMux I__2717 (
            .O(N__12440),
            .I(N__12421));
    LocalMux I__2716 (
            .O(N__12437),
            .I(N__12421));
    InMux I__2715 (
            .O(N__12436),
            .I(N__12418));
    LocalMux I__2714 (
            .O(N__12433),
            .I(N__12415));
    Span4Mux_h I__2713 (
            .O(N__12430),
            .I(N__12412));
    InMux I__2712 (
            .O(N__12429),
            .I(N__12409));
    Span4Mux_h I__2711 (
            .O(N__12426),
            .I(N__12404));
    Span4Mux_v I__2710 (
            .O(N__12421),
            .I(N__12404));
    LocalMux I__2709 (
            .O(N__12418),
            .I(N__12399));
    Span4Mux_v I__2708 (
            .O(N__12415),
            .I(N__12399));
    Odrv4 I__2707 (
            .O(N__12412),
            .I(ten_secsZ0Z_0));
    LocalMux I__2706 (
            .O(N__12409),
            .I(ten_secsZ0Z_0));
    Odrv4 I__2705 (
            .O(N__12404),
            .I(ten_secsZ0Z_0));
    Odrv4 I__2704 (
            .O(N__12399),
            .I(ten_secsZ0Z_0));
    CascadeMux I__2703 (
            .O(N__12390),
            .I(N__12387));
    InMux I__2702 (
            .O(N__12387),
            .I(N__12384));
    LocalMux I__2701 (
            .O(N__12384),
            .I(N__12381));
    Span4Mux_v I__2700 (
            .O(N__12381),
            .I(N__12378));
    Span4Mux_h I__2699 (
            .O(N__12378),
            .I(N__12375));
    Odrv4 I__2698 (
            .O(N__12375),
            .I(BNC1));
    InMux I__2697 (
            .O(N__12372),
            .I(N__12367));
    InMux I__2696 (
            .O(N__12371),
            .I(N__12362));
    InMux I__2695 (
            .O(N__12370),
            .I(N__12362));
    LocalMux I__2694 (
            .O(N__12367),
            .I(\d2.countZ0Z_9 ));
    LocalMux I__2693 (
            .O(N__12362),
            .I(\d2.countZ0Z_9 ));
    CascadeMux I__2692 (
            .O(N__12357),
            .I(N__12353));
    InMux I__2691 (
            .O(N__12356),
            .I(N__12349));
    InMux I__2690 (
            .O(N__12353),
            .I(N__12345));
    InMux I__2689 (
            .O(N__12352),
            .I(N__12342));
    LocalMux I__2688 (
            .O(N__12349),
            .I(N__12338));
    CascadeMux I__2687 (
            .O(N__12348),
            .I(N__12334));
    LocalMux I__2686 (
            .O(N__12345),
            .I(N__12331));
    LocalMux I__2685 (
            .O(N__12342),
            .I(N__12328));
    InMux I__2684 (
            .O(N__12341),
            .I(N__12323));
    Span4Mux_h I__2683 (
            .O(N__12338),
            .I(N__12320));
    InMux I__2682 (
            .O(N__12337),
            .I(N__12315));
    InMux I__2681 (
            .O(N__12334),
            .I(N__12315));
    Span4Mux_v I__2680 (
            .O(N__12331),
            .I(N__12310));
    Span4Mux_h I__2679 (
            .O(N__12328),
            .I(N__12310));
    InMux I__2678 (
            .O(N__12327),
            .I(N__12305));
    InMux I__2677 (
            .O(N__12326),
            .I(N__12305));
    LocalMux I__2676 (
            .O(N__12323),
            .I(d2_count_16));
    Odrv4 I__2675 (
            .O(N__12320),
            .I(d2_count_16));
    LocalMux I__2674 (
            .O(N__12315),
            .I(d2_count_16));
    Odrv4 I__2673 (
            .O(N__12310),
            .I(d2_count_16));
    LocalMux I__2672 (
            .O(N__12305),
            .I(d2_count_16));
    CascadeMux I__2671 (
            .O(N__12294),
            .I(N__12289));
    CascadeMux I__2670 (
            .O(N__12293),
            .I(N__12286));
    InMux I__2669 (
            .O(N__12292),
            .I(N__12283));
    InMux I__2668 (
            .O(N__12289),
            .I(N__12278));
    InMux I__2667 (
            .O(N__12286),
            .I(N__12278));
    LocalMux I__2666 (
            .O(N__12283),
            .I(\d2.countZ0Z_10 ));
    LocalMux I__2665 (
            .O(N__12278),
            .I(\d2.countZ0Z_10 ));
    InMux I__2664 (
            .O(N__12273),
            .I(N__12268));
    InMux I__2663 (
            .O(N__12272),
            .I(N__12263));
    InMux I__2662 (
            .O(N__12271),
            .I(N__12263));
    LocalMux I__2661 (
            .O(N__12268),
            .I(\d2.countZ0Z_7 ));
    LocalMux I__2660 (
            .O(N__12263),
            .I(\d2.countZ0Z_7 ));
    InMux I__2659 (
            .O(N__12258),
            .I(N__12255));
    LocalMux I__2658 (
            .O(N__12255),
            .I(N__12252));
    Odrv4 I__2657 (
            .O(N__12252),
            .I(\d2.g0_0_13 ));
    InMux I__2656 (
            .O(N__12249),
            .I(N__12239));
    InMux I__2655 (
            .O(N__12248),
            .I(N__12236));
    InMux I__2654 (
            .O(N__12247),
            .I(N__12233));
    InMux I__2653 (
            .O(N__12246),
            .I(N__12228));
    InMux I__2652 (
            .O(N__12245),
            .I(N__12228));
    InMux I__2651 (
            .O(N__12244),
            .I(N__12223));
    InMux I__2650 (
            .O(N__12243),
            .I(N__12223));
    InMux I__2649 (
            .O(N__12242),
            .I(N__12220));
    LocalMux I__2648 (
            .O(N__12239),
            .I(N__12217));
    LocalMux I__2647 (
            .O(N__12236),
            .I(d2_count_3));
    LocalMux I__2646 (
            .O(N__12233),
            .I(d2_count_3));
    LocalMux I__2645 (
            .O(N__12228),
            .I(d2_count_3));
    LocalMux I__2644 (
            .O(N__12223),
            .I(d2_count_3));
    LocalMux I__2643 (
            .O(N__12220),
            .I(d2_count_3));
    Odrv4 I__2642 (
            .O(N__12217),
            .I(d2_count_3));
    InMux I__2641 (
            .O(N__12204),
            .I(N__12201));
    LocalMux I__2640 (
            .O(N__12201),
            .I(\d1.g2_8_2 ));
    CascadeMux I__2639 (
            .O(N__12198),
            .I(N__12194));
    InMux I__2638 (
            .O(N__12197),
            .I(N__12190));
    InMux I__2637 (
            .O(N__12194),
            .I(N__12187));
    InMux I__2636 (
            .O(N__12193),
            .I(N__12184));
    LocalMux I__2635 (
            .O(N__12190),
            .I(\d2.countZ0Z_12 ));
    LocalMux I__2634 (
            .O(N__12187),
            .I(\d2.countZ0Z_12 ));
    LocalMux I__2633 (
            .O(N__12184),
            .I(\d2.countZ0Z_12 ));
    CascadeMux I__2632 (
            .O(N__12177),
            .I(N__12172));
    InMux I__2631 (
            .O(N__12176),
            .I(N__12169));
    InMux I__2630 (
            .O(N__12175),
            .I(N__12166));
    InMux I__2629 (
            .O(N__12172),
            .I(N__12163));
    LocalMux I__2628 (
            .O(N__12169),
            .I(\d2.countZ0Z_13 ));
    LocalMux I__2627 (
            .O(N__12166),
            .I(\d2.countZ0Z_13 ));
    LocalMux I__2626 (
            .O(N__12163),
            .I(\d2.countZ0Z_13 ));
    CascadeMux I__2625 (
            .O(N__12156),
            .I(N__12152));
    InMux I__2624 (
            .O(N__12155),
            .I(N__12148));
    InMux I__2623 (
            .O(N__12152),
            .I(N__12145));
    InMux I__2622 (
            .O(N__12151),
            .I(N__12142));
    LocalMux I__2621 (
            .O(N__12148),
            .I(\d2.countZ0Z_14 ));
    LocalMux I__2620 (
            .O(N__12145),
            .I(\d2.countZ0Z_14 ));
    LocalMux I__2619 (
            .O(N__12142),
            .I(\d2.countZ0Z_14 ));
    InMux I__2618 (
            .O(N__12135),
            .I(N__12131));
    InMux I__2617 (
            .O(N__12134),
            .I(N__12127));
    LocalMux I__2616 (
            .O(N__12131),
            .I(N__12124));
    InMux I__2615 (
            .O(N__12130),
            .I(N__12121));
    LocalMux I__2614 (
            .O(N__12127),
            .I(\d2.countZ0Z_11 ));
    Odrv4 I__2613 (
            .O(N__12124),
            .I(\d2.countZ0Z_11 ));
    LocalMux I__2612 (
            .O(N__12121),
            .I(\d2.countZ0Z_11 ));
    InMux I__2611 (
            .O(N__12114),
            .I(N__12110));
    InMux I__2610 (
            .O(N__12113),
            .I(N__12106));
    LocalMux I__2609 (
            .O(N__12110),
            .I(N__12103));
    InMux I__2608 (
            .O(N__12109),
            .I(N__12097));
    LocalMux I__2607 (
            .O(N__12106),
            .I(N__12093));
    Span4Mux_h I__2606 (
            .O(N__12103),
            .I(N__12090));
    CascadeMux I__2605 (
            .O(N__12102),
            .I(N__12087));
    InMux I__2604 (
            .O(N__12101),
            .I(N__12082));
    InMux I__2603 (
            .O(N__12100),
            .I(N__12082));
    LocalMux I__2602 (
            .O(N__12097),
            .I(N__12079));
    InMux I__2601 (
            .O(N__12096),
            .I(N__12076));
    Span4Mux_h I__2600 (
            .O(N__12093),
            .I(N__12071));
    Span4Mux_h I__2599 (
            .O(N__12090),
            .I(N__12071));
    InMux I__2598 (
            .O(N__12087),
            .I(N__12068));
    LocalMux I__2597 (
            .O(N__12082),
            .I(N__12063));
    Span4Mux_h I__2596 (
            .O(N__12079),
            .I(N__12063));
    LocalMux I__2595 (
            .O(N__12076),
            .I(d2_trans_up_1_15_7));
    Odrv4 I__2594 (
            .O(N__12071),
            .I(d2_trans_up_1_15_7));
    LocalMux I__2593 (
            .O(N__12068),
            .I(d2_trans_up_1_15_7));
    Odrv4 I__2592 (
            .O(N__12063),
            .I(d2_trans_up_1_15_7));
    InMux I__2591 (
            .O(N__12054),
            .I(N__12051));
    LocalMux I__2590 (
            .O(N__12051),
            .I(\d1.g2_i_a5_1Z0Z_6 ));
    InMux I__2589 (
            .O(N__12048),
            .I(N__12042));
    InMux I__2588 (
            .O(N__12047),
            .I(N__12039));
    CascadeMux I__2587 (
            .O(N__12046),
            .I(N__12036));
    CascadeMux I__2586 (
            .O(N__12045),
            .I(N__12033));
    LocalMux I__2585 (
            .O(N__12042),
            .I(N__12029));
    LocalMux I__2584 (
            .O(N__12039),
            .I(N__12026));
    InMux I__2583 (
            .O(N__12036),
            .I(N__12022));
    InMux I__2582 (
            .O(N__12033),
            .I(N__12019));
    CascadeMux I__2581 (
            .O(N__12032),
            .I(N__12014));
    Span4Mux_h I__2580 (
            .O(N__12029),
            .I(N__12009));
    Span4Mux_h I__2579 (
            .O(N__12026),
            .I(N__12009));
    InMux I__2578 (
            .O(N__12025),
            .I(N__12006));
    LocalMux I__2577 (
            .O(N__12022),
            .I(N__12001));
    LocalMux I__2576 (
            .O(N__12019),
            .I(N__12001));
    InMux I__2575 (
            .O(N__12018),
            .I(N__11994));
    InMux I__2574 (
            .O(N__12017),
            .I(N__11994));
    InMux I__2573 (
            .O(N__12014),
            .I(N__11994));
    Odrv4 I__2572 (
            .O(N__12009),
            .I(d2_sync_1));
    LocalMux I__2571 (
            .O(N__12006),
            .I(d2_sync_1));
    Odrv12 I__2570 (
            .O(N__12001),
            .I(d2_sync_1));
    LocalMux I__2569 (
            .O(N__11994),
            .I(d2_sync_1));
    CascadeMux I__2568 (
            .O(N__11985),
            .I(N__11982));
    InMux I__2567 (
            .O(N__11982),
            .I(N__11977));
    InMux I__2566 (
            .O(N__11981),
            .I(N__11974));
    InMux I__2565 (
            .O(N__11980),
            .I(N__11969));
    LocalMux I__2564 (
            .O(N__11977),
            .I(N__11964));
    LocalMux I__2563 (
            .O(N__11974),
            .I(N__11964));
    InMux I__2562 (
            .O(N__11973),
            .I(N__11959));
    InMux I__2561 (
            .O(N__11972),
            .I(N__11959));
    LocalMux I__2560 (
            .O(N__11969),
            .I(N__11955));
    Span4Mux_v I__2559 (
            .O(N__11964),
            .I(N__11950));
    LocalMux I__2558 (
            .O(N__11959),
            .I(N__11950));
    CascadeMux I__2557 (
            .O(N__11958),
            .I(N__11946));
    Span4Mux_v I__2556 (
            .O(N__11955),
            .I(N__11940));
    Span4Mux_h I__2555 (
            .O(N__11950),
            .I(N__11940));
    InMux I__2554 (
            .O(N__11949),
            .I(N__11933));
    InMux I__2553 (
            .O(N__11946),
            .I(N__11933));
    InMux I__2552 (
            .O(N__11945),
            .I(N__11933));
    Odrv4 I__2551 (
            .O(N__11940),
            .I(d2_state));
    LocalMux I__2550 (
            .O(N__11933),
            .I(d2_state));
    IoInMux I__2549 (
            .O(N__11928),
            .I(N__11925));
    LocalMux I__2548 (
            .O(N__11925),
            .I(N__11922));
    Odrv12 I__2547 (
            .O(N__11922),
            .I(\d2.idle_i ));
    InMux I__2546 (
            .O(N__11919),
            .I(N__11915));
    InMux I__2545 (
            .O(N__11918),
            .I(N__11912));
    LocalMux I__2544 (
            .O(N__11915),
            .I(d2_g0_3));
    LocalMux I__2543 (
            .O(N__11912),
            .I(d2_g0_3));
    CascadeMux I__2542 (
            .O(N__11907),
            .I(\d1.g0_1_0_a4Z0Z_4_cascade_ ));
    InMux I__2541 (
            .O(N__11904),
            .I(N__11895));
    InMux I__2540 (
            .O(N__11903),
            .I(N__11892));
    InMux I__2539 (
            .O(N__11902),
            .I(N__11883));
    InMux I__2538 (
            .O(N__11901),
            .I(N__11878));
    InMux I__2537 (
            .O(N__11900),
            .I(N__11873));
    InMux I__2536 (
            .O(N__11899),
            .I(N__11873));
    InMux I__2535 (
            .O(N__11898),
            .I(N__11870));
    LocalMux I__2534 (
            .O(N__11895),
            .I(N__11865));
    LocalMux I__2533 (
            .O(N__11892),
            .I(N__11865));
    InMux I__2532 (
            .O(N__11891),
            .I(N__11853));
    InMux I__2531 (
            .O(N__11890),
            .I(N__11853));
    InMux I__2530 (
            .O(N__11889),
            .I(N__11853));
    InMux I__2529 (
            .O(N__11888),
            .I(N__11846));
    InMux I__2528 (
            .O(N__11887),
            .I(N__11846));
    InMux I__2527 (
            .O(N__11886),
            .I(N__11846));
    LocalMux I__2526 (
            .O(N__11883),
            .I(N__11843));
    InMux I__2525 (
            .O(N__11882),
            .I(N__11838));
    InMux I__2524 (
            .O(N__11881),
            .I(N__11838));
    LocalMux I__2523 (
            .O(N__11878),
            .I(N__11829));
    LocalMux I__2522 (
            .O(N__11873),
            .I(N__11829));
    LocalMux I__2521 (
            .O(N__11870),
            .I(N__11829));
    Span4Mux_h I__2520 (
            .O(N__11865),
            .I(N__11829));
    InMux I__2519 (
            .O(N__11864),
            .I(N__11826));
    InMux I__2518 (
            .O(N__11863),
            .I(N__11823));
    InMux I__2517 (
            .O(N__11862),
            .I(N__11818));
    InMux I__2516 (
            .O(N__11861),
            .I(N__11818));
    InMux I__2515 (
            .O(N__11860),
            .I(N__11815));
    LocalMux I__2514 (
            .O(N__11853),
            .I(N__11810));
    LocalMux I__2513 (
            .O(N__11846),
            .I(N__11810));
    Span4Mux_v I__2512 (
            .O(N__11843),
            .I(N__11807));
    LocalMux I__2511 (
            .O(N__11838),
            .I(N__11804));
    Span4Mux_v I__2510 (
            .O(N__11829),
            .I(N__11801));
    LocalMux I__2509 (
            .O(N__11826),
            .I(N__11794));
    LocalMux I__2508 (
            .O(N__11823),
            .I(N__11794));
    LocalMux I__2507 (
            .O(N__11818),
            .I(N__11794));
    LocalMux I__2506 (
            .O(N__11815),
            .I(N__11791));
    Span4Mux_v I__2505 (
            .O(N__11810),
            .I(N__11784));
    Span4Mux_h I__2504 (
            .O(N__11807),
            .I(N__11784));
    Span4Mux_v I__2503 (
            .O(N__11804),
            .I(N__11784));
    Odrv4 I__2502 (
            .O(N__11801),
            .I(stateZ0Z_1));
    Odrv12 I__2501 (
            .O(N__11794),
            .I(stateZ0Z_1));
    Odrv4 I__2500 (
            .O(N__11791),
            .I(stateZ0Z_1));
    Odrv4 I__2499 (
            .O(N__11784),
            .I(stateZ0Z_1));
    InMux I__2498 (
            .O(N__11775),
            .I(N__11772));
    LocalMux I__2497 (
            .O(N__11772),
            .I(N__11769));
    Odrv12 I__2496 (
            .O(N__11769),
            .I(\d1.g0_1_0_a4Z0Z_8 ));
    CascadeMux I__2495 (
            .O(N__11766),
            .I(N__11762));
    InMux I__2494 (
            .O(N__11765),
            .I(N__11754));
    InMux I__2493 (
            .O(N__11762),
            .I(N__11754));
    CascadeMux I__2492 (
            .O(N__11761),
            .I(N__11748));
    InMux I__2491 (
            .O(N__11760),
            .I(N__11744));
    InMux I__2490 (
            .O(N__11759),
            .I(N__11741));
    LocalMux I__2489 (
            .O(N__11754),
            .I(N__11738));
    InMux I__2488 (
            .O(N__11753),
            .I(N__11735));
    InMux I__2487 (
            .O(N__11752),
            .I(N__11728));
    InMux I__2486 (
            .O(N__11751),
            .I(N__11728));
    InMux I__2485 (
            .O(N__11748),
            .I(N__11728));
    InMux I__2484 (
            .O(N__11747),
            .I(N__11725));
    LocalMux I__2483 (
            .O(N__11744),
            .I(d2_count_15));
    LocalMux I__2482 (
            .O(N__11741),
            .I(d2_count_15));
    Odrv4 I__2481 (
            .O(N__11738),
            .I(d2_count_15));
    LocalMux I__2480 (
            .O(N__11735),
            .I(d2_count_15));
    LocalMux I__2479 (
            .O(N__11728),
            .I(d2_count_15));
    LocalMux I__2478 (
            .O(N__11725),
            .I(d2_count_15));
    CascadeMux I__2477 (
            .O(N__11712),
            .I(N__11707));
    CascadeMux I__2476 (
            .O(N__11711),
            .I(N__11704));
    InMux I__2475 (
            .O(N__11710),
            .I(N__11701));
    InMux I__2474 (
            .O(N__11707),
            .I(N__11698));
    InMux I__2473 (
            .O(N__11704),
            .I(N__11691));
    LocalMux I__2472 (
            .O(N__11701),
            .I(N__11686));
    LocalMux I__2471 (
            .O(N__11698),
            .I(N__11686));
    CascadeMux I__2470 (
            .O(N__11697),
            .I(N__11681));
    InMux I__2469 (
            .O(N__11696),
            .I(N__11677));
    InMux I__2468 (
            .O(N__11695),
            .I(N__11674));
    InMux I__2467 (
            .O(N__11694),
            .I(N__11671));
    LocalMux I__2466 (
            .O(N__11691),
            .I(N__11666));
    Span4Mux_v I__2465 (
            .O(N__11686),
            .I(N__11666));
    InMux I__2464 (
            .O(N__11685),
            .I(N__11661));
    InMux I__2463 (
            .O(N__11684),
            .I(N__11661));
    InMux I__2462 (
            .O(N__11681),
            .I(N__11656));
    InMux I__2461 (
            .O(N__11680),
            .I(N__11656));
    LocalMux I__2460 (
            .O(N__11677),
            .I(d2_count_2));
    LocalMux I__2459 (
            .O(N__11674),
            .I(d2_count_2));
    LocalMux I__2458 (
            .O(N__11671),
            .I(d2_count_2));
    Odrv4 I__2457 (
            .O(N__11666),
            .I(d2_count_2));
    LocalMux I__2456 (
            .O(N__11661),
            .I(d2_count_2));
    LocalMux I__2455 (
            .O(N__11656),
            .I(d2_count_2));
    CascadeMux I__2454 (
            .O(N__11643),
            .I(N__11640));
    InMux I__2453 (
            .O(N__11640),
            .I(N__11635));
    InMux I__2452 (
            .O(N__11639),
            .I(N__11629));
    InMux I__2451 (
            .O(N__11638),
            .I(N__11629));
    LocalMux I__2450 (
            .O(N__11635),
            .I(N__11623));
    InMux I__2449 (
            .O(N__11634),
            .I(N__11617));
    LocalMux I__2448 (
            .O(N__11629),
            .I(N__11614));
    InMux I__2447 (
            .O(N__11628),
            .I(N__11609));
    InMux I__2446 (
            .O(N__11627),
            .I(N__11609));
    InMux I__2445 (
            .O(N__11626),
            .I(N__11605));
    Span4Mux_h I__2444 (
            .O(N__11623),
            .I(N__11602));
    InMux I__2443 (
            .O(N__11622),
            .I(N__11599));
    InMux I__2442 (
            .O(N__11621),
            .I(N__11594));
    InMux I__2441 (
            .O(N__11620),
            .I(N__11594));
    LocalMux I__2440 (
            .O(N__11617),
            .I(N__11591));
    Span4Mux_v I__2439 (
            .O(N__11614),
            .I(N__11586));
    LocalMux I__2438 (
            .O(N__11609),
            .I(N__11586));
    InMux I__2437 (
            .O(N__11608),
            .I(N__11583));
    LocalMux I__2436 (
            .O(N__11605),
            .I(d2_count_1));
    Odrv4 I__2435 (
            .O(N__11602),
            .I(d2_count_1));
    LocalMux I__2434 (
            .O(N__11599),
            .I(d2_count_1));
    LocalMux I__2433 (
            .O(N__11594),
            .I(d2_count_1));
    Odrv4 I__2432 (
            .O(N__11591),
            .I(d2_count_1));
    Odrv4 I__2431 (
            .O(N__11586),
            .I(d2_count_1));
    LocalMux I__2430 (
            .O(N__11583),
            .I(d2_count_1));
    SRMux I__2429 (
            .O(N__11568),
            .I(N__11565));
    LocalMux I__2428 (
            .O(N__11565),
            .I(N__11561));
    SRMux I__2427 (
            .O(N__11564),
            .I(N__11558));
    Span4Mux_h I__2426 (
            .O(N__11561),
            .I(N__11555));
    LocalMux I__2425 (
            .O(N__11558),
            .I(N__11552));
    Span4Mux_h I__2424 (
            .O(N__11555),
            .I(N__11548));
    Span4Mux_v I__2423 (
            .O(N__11552),
            .I(N__11545));
    SRMux I__2422 (
            .O(N__11551),
            .I(N__11542));
    Span4Mux_h I__2421 (
            .O(N__11548),
            .I(N__11538));
    Span4Mux_h I__2420 (
            .O(N__11545),
            .I(N__11535));
    LocalMux I__2419 (
            .O(N__11542),
            .I(N__11532));
    InMux I__2418 (
            .O(N__11541),
            .I(N__11529));
    Odrv4 I__2417 (
            .O(N__11538),
            .I(mins_0_sqmuxa));
    Odrv4 I__2416 (
            .O(N__11535),
            .I(mins_0_sqmuxa));
    Odrv12 I__2415 (
            .O(N__11532),
            .I(mins_0_sqmuxa));
    LocalMux I__2414 (
            .O(N__11529),
            .I(mins_0_sqmuxa));
    CascadeMux I__2413 (
            .O(N__11520),
            .I(N__11517));
    InMux I__2412 (
            .O(N__11517),
            .I(N__11514));
    LocalMux I__2411 (
            .O(N__11514),
            .I(N__11511));
    Span4Mux_h I__2410 (
            .O(N__11511),
            .I(N__11508));
    Odrv4 I__2409 (
            .O(N__11508),
            .I(\d1.g0_1_a5_0Z0Z_11 ));
    InMux I__2408 (
            .O(N__11505),
            .I(N__11502));
    LocalMux I__2407 (
            .O(N__11502),
            .I(N__11499));
    Span4Mux_v I__2406 (
            .O(N__11499),
            .I(N__11496));
    Odrv4 I__2405 (
            .O(N__11496),
            .I(\d1.g2_12_1 ));
    InMux I__2404 (
            .O(N__11493),
            .I(N__11489));
    InMux I__2403 (
            .O(N__11492),
            .I(N__11485));
    LocalMux I__2402 (
            .O(N__11489),
            .I(N__11481));
    InMux I__2401 (
            .O(N__11488),
            .I(N__11475));
    LocalMux I__2400 (
            .O(N__11485),
            .I(N__11472));
    InMux I__2399 (
            .O(N__11484),
            .I(N__11469));
    Span4Mux_h I__2398 (
            .O(N__11481),
            .I(N__11466));
    InMux I__2397 (
            .O(N__11480),
            .I(N__11459));
    InMux I__2396 (
            .O(N__11479),
            .I(N__11459));
    InMux I__2395 (
            .O(N__11478),
            .I(N__11459));
    LocalMux I__2394 (
            .O(N__11475),
            .I(d2_count_4));
    Odrv4 I__2393 (
            .O(N__11472),
            .I(d2_count_4));
    LocalMux I__2392 (
            .O(N__11469),
            .I(d2_count_4));
    Odrv4 I__2391 (
            .O(N__11466),
            .I(d2_count_4));
    LocalMux I__2390 (
            .O(N__11459),
            .I(d2_count_4));
    InMux I__2389 (
            .O(N__11448),
            .I(N__11444));
    InMux I__2388 (
            .O(N__11447),
            .I(N__11441));
    LocalMux I__2387 (
            .O(N__11444),
            .I(N__11435));
    LocalMux I__2386 (
            .O(N__11441),
            .I(N__11431));
    InMux I__2385 (
            .O(N__11440),
            .I(N__11428));
    InMux I__2384 (
            .O(N__11439),
            .I(N__11420));
    InMux I__2383 (
            .O(N__11438),
            .I(N__11420));
    Span4Mux_h I__2382 (
            .O(N__11435),
            .I(N__11417));
    InMux I__2381 (
            .O(N__11434),
            .I(N__11414));
    Span4Mux_h I__2380 (
            .O(N__11431),
            .I(N__11411));
    LocalMux I__2379 (
            .O(N__11428),
            .I(N__11408));
    InMux I__2378 (
            .O(N__11427),
            .I(N__11401));
    InMux I__2377 (
            .O(N__11426),
            .I(N__11401));
    InMux I__2376 (
            .O(N__11425),
            .I(N__11401));
    LocalMux I__2375 (
            .O(N__11420),
            .I(d2_count_0));
    Odrv4 I__2374 (
            .O(N__11417),
            .I(d2_count_0));
    LocalMux I__2373 (
            .O(N__11414),
            .I(d2_count_0));
    Odrv4 I__2372 (
            .O(N__11411),
            .I(d2_count_0));
    Odrv4 I__2371 (
            .O(N__11408),
            .I(d2_count_0));
    LocalMux I__2370 (
            .O(N__11401),
            .I(d2_count_0));
    InMux I__2369 (
            .O(N__11388),
            .I(N__11385));
    LocalMux I__2368 (
            .O(N__11385),
            .I(N__11382));
    Span4Mux_v I__2367 (
            .O(N__11382),
            .I(N__11379));
    Span4Mux_h I__2366 (
            .O(N__11379),
            .I(N__11376));
    Odrv4 I__2365 (
            .O(N__11376),
            .I(\d2.trans_up_1_15 ));
    CascadeMux I__2364 (
            .O(N__11373),
            .I(\d2.trans_up_1_15_cascade_ ));
    InMux I__2363 (
            .O(N__11370),
            .I(N__11367));
    LocalMux I__2362 (
            .O(N__11367),
            .I(s_dn_0));
    InMux I__2361 (
            .O(N__11364),
            .I(N__11361));
    LocalMux I__2360 (
            .O(N__11361),
            .I(\d1.g2Z0Z_8 ));
    CascadeMux I__2359 (
            .O(N__11358),
            .I(N__11355));
    InMux I__2358 (
            .O(N__11355),
            .I(N__11352));
    LocalMux I__2357 (
            .O(N__11352),
            .I(\d1.mins27_0_0 ));
    InMux I__2356 (
            .O(N__11349),
            .I(N__11346));
    LocalMux I__2355 (
            .O(N__11346),
            .I(\d1.g2_i_a5_0Z0Z_7 ));
    InMux I__2354 (
            .O(N__11343),
            .I(N__11339));
    InMux I__2353 (
            .O(N__11342),
            .I(N__11336));
    LocalMux I__2352 (
            .O(N__11339),
            .I(N__11332));
    LocalMux I__2351 (
            .O(N__11336),
            .I(N__11329));
    InMux I__2350 (
            .O(N__11335),
            .I(N__11326));
    Span4Mux_h I__2349 (
            .O(N__11332),
            .I(N__11323));
    Odrv12 I__2348 (
            .O(N__11329),
            .I(d2_trans_up_1_15_1));
    LocalMux I__2347 (
            .O(N__11326),
            .I(d2_trans_up_1_15_1));
    Odrv4 I__2346 (
            .O(N__11323),
            .I(d2_trans_up_1_15_1));
    CascadeMux I__2345 (
            .O(N__11316),
            .I(d2_g0_3_cascade_));
    InMux I__2344 (
            .O(N__11313),
            .I(N__11310));
    LocalMux I__2343 (
            .O(N__11310),
            .I(\d1.g2_i_a5_1Z0Z_7 ));
    InMux I__2342 (
            .O(N__11307),
            .I(N__11303));
    InMux I__2341 (
            .O(N__11306),
            .I(N__11300));
    LocalMux I__2340 (
            .O(N__11303),
            .I(N__11294));
    LocalMux I__2339 (
            .O(N__11300),
            .I(N__11294));
    InMux I__2338 (
            .O(N__11299),
            .I(N__11291));
    Odrv4 I__2337 (
            .O(N__11294),
            .I(\d2.countZ0Z_8 ));
    LocalMux I__2336 (
            .O(N__11291),
            .I(\d2.countZ0Z_8 ));
    InMux I__2335 (
            .O(N__11286),
            .I(N__11281));
    InMux I__2334 (
            .O(N__11285),
            .I(N__11276));
    InMux I__2333 (
            .O(N__11284),
            .I(N__11276));
    LocalMux I__2332 (
            .O(N__11281),
            .I(N__11273));
    LocalMux I__2331 (
            .O(N__11276),
            .I(N__11266));
    Span4Mux_h I__2330 (
            .O(N__11273),
            .I(N__11263));
    InMux I__2329 (
            .O(N__11272),
            .I(N__11260));
    InMux I__2328 (
            .O(N__11271),
            .I(N__11255));
    InMux I__2327 (
            .O(N__11270),
            .I(N__11255));
    InMux I__2326 (
            .O(N__11269),
            .I(N__11252));
    Span4Mux_v I__2325 (
            .O(N__11266),
            .I(N__11249));
    Odrv4 I__2324 (
            .O(N__11263),
            .I(d2_trans_up_1_15_8));
    LocalMux I__2323 (
            .O(N__11260),
            .I(d2_trans_up_1_15_8));
    LocalMux I__2322 (
            .O(N__11255),
            .I(d2_trans_up_1_15_8));
    LocalMux I__2321 (
            .O(N__11252),
            .I(d2_trans_up_1_15_8));
    Odrv4 I__2320 (
            .O(N__11249),
            .I(d2_trans_up_1_15_8));
    InMux I__2319 (
            .O(N__11238),
            .I(N__11234));
    InMux I__2318 (
            .O(N__11237),
            .I(N__11231));
    LocalMux I__2317 (
            .O(N__11234),
            .I(N__11225));
    LocalMux I__2316 (
            .O(N__11231),
            .I(N__11222));
    CascadeMux I__2315 (
            .O(N__11230),
            .I(N__11218));
    InMux I__2314 (
            .O(N__11229),
            .I(N__11214));
    InMux I__2313 (
            .O(N__11228),
            .I(N__11211));
    Span4Mux_v I__2312 (
            .O(N__11225),
            .I(N__11208));
    Span4Mux_h I__2311 (
            .O(N__11222),
            .I(N__11205));
    InMux I__2310 (
            .O(N__11221),
            .I(N__11200));
    InMux I__2309 (
            .O(N__11218),
            .I(N__11200));
    InMux I__2308 (
            .O(N__11217),
            .I(N__11197));
    LocalMux I__2307 (
            .O(N__11214),
            .I(N__11194));
    LocalMux I__2306 (
            .O(N__11211),
            .I(d2_count_6));
    Odrv4 I__2305 (
            .O(N__11208),
            .I(d2_count_6));
    Odrv4 I__2304 (
            .O(N__11205),
            .I(d2_count_6));
    LocalMux I__2303 (
            .O(N__11200),
            .I(d2_count_6));
    LocalMux I__2302 (
            .O(N__11197),
            .I(d2_count_6));
    Odrv4 I__2301 (
            .O(N__11194),
            .I(d2_count_6));
    InMux I__2300 (
            .O(N__11181),
            .I(N__11177));
    InMux I__2299 (
            .O(N__11180),
            .I(N__11174));
    LocalMux I__2298 (
            .O(N__11177),
            .I(N__11169));
    LocalMux I__2297 (
            .O(N__11174),
            .I(N__11166));
    InMux I__2296 (
            .O(N__11173),
            .I(N__11160));
    InMux I__2295 (
            .O(N__11172),
            .I(N__11157));
    Span4Mux_v I__2294 (
            .O(N__11169),
            .I(N__11154));
    Span4Mux_h I__2293 (
            .O(N__11166),
            .I(N__11151));
    InMux I__2292 (
            .O(N__11165),
            .I(N__11146));
    InMux I__2291 (
            .O(N__11164),
            .I(N__11146));
    InMux I__2290 (
            .O(N__11163),
            .I(N__11143));
    LocalMux I__2289 (
            .O(N__11160),
            .I(N__11140));
    LocalMux I__2288 (
            .O(N__11157),
            .I(d2_count_5));
    Odrv4 I__2287 (
            .O(N__11154),
            .I(d2_count_5));
    Odrv4 I__2286 (
            .O(N__11151),
            .I(d2_count_5));
    LocalMux I__2285 (
            .O(N__11146),
            .I(d2_count_5));
    LocalMux I__2284 (
            .O(N__11143),
            .I(d2_count_5));
    Odrv4 I__2283 (
            .O(N__11140),
            .I(d2_count_5));
    CascadeMux I__2282 (
            .O(N__11127),
            .I(\d1.g2_7_0_cascade_ ));
    InMux I__2281 (
            .O(N__11124),
            .I(N__11121));
    LocalMux I__2280 (
            .O(N__11121),
            .I(N__11118));
    Odrv12 I__2279 (
            .O(N__11118),
            .I(\d1.g2_11_0 ));
    InMux I__2278 (
            .O(N__11115),
            .I(N__11112));
    LocalMux I__2277 (
            .O(N__11112),
            .I(N__11109));
    Odrv12 I__2276 (
            .O(N__11109),
            .I(\d1.N_3 ));
    CascadeMux I__2275 (
            .O(N__11106),
            .I(N__11103));
    InMux I__2274 (
            .O(N__11103),
            .I(N__11100));
    LocalMux I__2273 (
            .O(N__11100),
            .I(N__11097));
    Span4Mux_h I__2272 (
            .O(N__11097),
            .I(N__11094));
    Odrv4 I__2271 (
            .O(N__11094),
            .I(\d3.trans_up_1_14_2 ));
    InMux I__2270 (
            .O(N__11091),
            .I(N__11088));
    LocalMux I__2269 (
            .O(N__11088),
            .I(N__11085));
    Span4Mux_h I__2268 (
            .O(N__11085),
            .I(N__11079));
    InMux I__2267 (
            .O(N__11084),
            .I(N__11076));
    InMux I__2266 (
            .O(N__11083),
            .I(N__11073));
    InMux I__2265 (
            .O(N__11082),
            .I(N__11070));
    Odrv4 I__2264 (
            .O(N__11079),
            .I(d3_trans_up_1_15));
    LocalMux I__2263 (
            .O(N__11076),
            .I(d3_trans_up_1_15));
    LocalMux I__2262 (
            .O(N__11073),
            .I(d3_trans_up_1_15));
    LocalMux I__2261 (
            .O(N__11070),
            .I(d3_trans_up_1_15));
    InMux I__2260 (
            .O(N__11061),
            .I(N__11058));
    LocalMux I__2259 (
            .O(N__11058),
            .I(N__11054));
    InMux I__2258 (
            .O(N__11057),
            .I(N__11049));
    Span4Mux_h I__2257 (
            .O(N__11054),
            .I(N__11046));
    InMux I__2256 (
            .O(N__11053),
            .I(N__11041));
    InMux I__2255 (
            .O(N__11052),
            .I(N__11041));
    LocalMux I__2254 (
            .O(N__11049),
            .I(\d1.countZ0Z_5 ));
    Odrv4 I__2253 (
            .O(N__11046),
            .I(\d1.countZ0Z_5 ));
    LocalMux I__2252 (
            .O(N__11041),
            .I(\d1.countZ0Z_5 ));
    InMux I__2251 (
            .O(N__11034),
            .I(N__11031));
    LocalMux I__2250 (
            .O(N__11031),
            .I(N__11027));
    InMux I__2249 (
            .O(N__11030),
            .I(N__11022));
    Span4Mux_h I__2248 (
            .O(N__11027),
            .I(N__11019));
    InMux I__2247 (
            .O(N__11026),
            .I(N__11014));
    InMux I__2246 (
            .O(N__11025),
            .I(N__11014));
    LocalMux I__2245 (
            .O(N__11022),
            .I(\d1.countZ0Z_4 ));
    Odrv4 I__2244 (
            .O(N__11019),
            .I(\d1.countZ0Z_4 ));
    LocalMux I__2243 (
            .O(N__11014),
            .I(\d1.countZ0Z_4 ));
    CascadeMux I__2242 (
            .O(N__11007),
            .I(N__11003));
    InMux I__2241 (
            .O(N__11006),
            .I(N__10998));
    InMux I__2240 (
            .O(N__11003),
            .I(N__10995));
    CascadeMux I__2239 (
            .O(N__11002),
            .I(N__10992));
    CascadeMux I__2238 (
            .O(N__11001),
            .I(N__10989));
    LocalMux I__2237 (
            .O(N__10998),
            .I(N__10984));
    LocalMux I__2236 (
            .O(N__10995),
            .I(N__10984));
    InMux I__2235 (
            .O(N__10992),
            .I(N__10979));
    InMux I__2234 (
            .O(N__10989),
            .I(N__10979));
    Odrv12 I__2233 (
            .O(N__10984),
            .I(\d1.countZ0Z_6 ));
    LocalMux I__2232 (
            .O(N__10979),
            .I(\d1.countZ0Z_6 ));
    InMux I__2231 (
            .O(N__10974),
            .I(N__10970));
    InMux I__2230 (
            .O(N__10973),
            .I(N__10965));
    LocalMux I__2229 (
            .O(N__10970),
            .I(N__10962));
    InMux I__2228 (
            .O(N__10969),
            .I(N__10957));
    InMux I__2227 (
            .O(N__10968),
            .I(N__10957));
    LocalMux I__2226 (
            .O(N__10965),
            .I(\d1.countZ0Z_3 ));
    Odrv12 I__2225 (
            .O(N__10962),
            .I(\d1.countZ0Z_3 ));
    LocalMux I__2224 (
            .O(N__10957),
            .I(\d1.countZ0Z_3 ));
    InMux I__2223 (
            .O(N__10950),
            .I(N__10947));
    LocalMux I__2222 (
            .O(N__10947),
            .I(N__10942));
    InMux I__2221 (
            .O(N__10946),
            .I(N__10939));
    CascadeMux I__2220 (
            .O(N__10945),
            .I(N__10936));
    Span4Mux_v I__2219 (
            .O(N__10942),
            .I(N__10933));
    LocalMux I__2218 (
            .O(N__10939),
            .I(N__10930));
    InMux I__2217 (
            .O(N__10936),
            .I(N__10927));
    Span4Mux_h I__2216 (
            .O(N__10933),
            .I(N__10924));
    Span4Mux_v I__2215 (
            .O(N__10930),
            .I(N__10919));
    LocalMux I__2214 (
            .O(N__10927),
            .I(N__10919));
    Odrv4 I__2213 (
            .O(N__10924),
            .I(\d1.trans_up_1_12 ));
    Odrv4 I__2212 (
            .O(N__10919),
            .I(\d1.trans_up_1_12 ));
    CascadeMux I__2211 (
            .O(N__10914),
            .I(\d1.g1_9_cascade_ ));
    InMux I__2210 (
            .O(N__10911),
            .I(N__10908));
    LocalMux I__2209 (
            .O(N__10908),
            .I(N__10905));
    Odrv12 I__2208 (
            .O(N__10905),
            .I(\d1.g1_13 ));
    InMux I__2207 (
            .O(N__10902),
            .I(N__10898));
    InMux I__2206 (
            .O(N__10901),
            .I(N__10893));
    LocalMux I__2205 (
            .O(N__10898),
            .I(N__10889));
    InMux I__2204 (
            .O(N__10897),
            .I(N__10886));
    InMux I__2203 (
            .O(N__10896),
            .I(N__10882));
    LocalMux I__2202 (
            .O(N__10893),
            .I(N__10879));
    InMux I__2201 (
            .O(N__10892),
            .I(N__10875));
    Span4Mux_h I__2200 (
            .O(N__10889),
            .I(N__10872));
    LocalMux I__2199 (
            .O(N__10886),
            .I(N__10869));
    InMux I__2198 (
            .O(N__10885),
            .I(N__10866));
    LocalMux I__2197 (
            .O(N__10882),
            .I(N__10861));
    Span4Mux_v I__2196 (
            .O(N__10879),
            .I(N__10861));
    InMux I__2195 (
            .O(N__10878),
            .I(N__10858));
    LocalMux I__2194 (
            .O(N__10875),
            .I(un1_alarm_on_0_sqmuxa_0));
    Odrv4 I__2193 (
            .O(N__10872),
            .I(un1_alarm_on_0_sqmuxa_0));
    Odrv4 I__2192 (
            .O(N__10869),
            .I(un1_alarm_on_0_sqmuxa_0));
    LocalMux I__2191 (
            .O(N__10866),
            .I(un1_alarm_on_0_sqmuxa_0));
    Odrv4 I__2190 (
            .O(N__10861),
            .I(un1_alarm_on_0_sqmuxa_0));
    LocalMux I__2189 (
            .O(N__10858),
            .I(un1_alarm_on_0_sqmuxa_0));
    InMux I__2188 (
            .O(N__10845),
            .I(N__10842));
    LocalMux I__2187 (
            .O(N__10842),
            .I(\d1.g2_iZ0Z_0 ));
    CascadeMux I__2186 (
            .O(N__10839),
            .I(N__10836));
    InMux I__2185 (
            .O(N__10836),
            .I(N__10833));
    LocalMux I__2184 (
            .O(N__10833),
            .I(\d1.N_6 ));
    InMux I__2183 (
            .O(N__10830),
            .I(N__10827));
    LocalMux I__2182 (
            .O(N__10827),
            .I(N__10822));
    CascadeMux I__2181 (
            .O(N__10826),
            .I(N__10819));
    InMux I__2180 (
            .O(N__10825),
            .I(N__10816));
    Span4Mux_h I__2179 (
            .O(N__10822),
            .I(N__10813));
    InMux I__2178 (
            .O(N__10819),
            .I(N__10810));
    LocalMux I__2177 (
            .O(N__10816),
            .I(ten_secs_1_sqmuxa));
    Odrv4 I__2176 (
            .O(N__10813),
            .I(ten_secs_1_sqmuxa));
    LocalMux I__2175 (
            .O(N__10810),
            .I(ten_secs_1_sqmuxa));
    InMux I__2174 (
            .O(N__10803),
            .I(N__10800));
    LocalMux I__2173 (
            .O(N__10800),
            .I(\d1.mins_2_sqmuxa_1 ));
    InMux I__2172 (
            .O(N__10797),
            .I(N__10794));
    LocalMux I__2171 (
            .O(N__10794),
            .I(\d1.mins_16_1Z0Z_3 ));
    CascadeMux I__2170 (
            .O(N__10791),
            .I(\d1.g3_0_cascade_ ));
    InMux I__2169 (
            .O(N__10788),
            .I(N__10785));
    LocalMux I__2168 (
            .O(N__10785),
            .I(\d1.N_8_0 ));
    CascadeMux I__2167 (
            .O(N__10782),
            .I(un1_state_0_sqmuxa_1_0_cascade_));
    SRMux I__2166 (
            .O(N__10779),
            .I(N__10775));
    CEMux I__2165 (
            .O(N__10778),
            .I(N__10771));
    LocalMux I__2164 (
            .O(N__10775),
            .I(N__10768));
    CEMux I__2163 (
            .O(N__10774),
            .I(N__10765));
    LocalMux I__2162 (
            .O(N__10771),
            .I(N__10762));
    Span4Mux_h I__2161 (
            .O(N__10768),
            .I(N__10759));
    LocalMux I__2160 (
            .O(N__10765),
            .I(N__10756));
    Span4Mux_h I__2159 (
            .O(N__10762),
            .I(N__10753));
    Span4Mux_h I__2158 (
            .O(N__10759),
            .I(N__10750));
    Odrv12 I__2157 (
            .O(N__10756),
            .I(mins_stored_0_sqmuxa));
    Odrv4 I__2156 (
            .O(N__10753),
            .I(mins_stored_0_sqmuxa));
    Odrv4 I__2155 (
            .O(N__10750),
            .I(mins_stored_0_sqmuxa));
    CascadeMux I__2154 (
            .O(N__10743),
            .I(N__10740));
    InMux I__2153 (
            .O(N__10740),
            .I(N__10737));
    LocalMux I__2152 (
            .O(N__10737),
            .I(N__10734));
    Odrv4 I__2151 (
            .O(N__10734),
            .I(\d1.state_0_sqmuxaZ0Z_1 ));
    InMux I__2150 (
            .O(N__10731),
            .I(N__10728));
    LocalMux I__2149 (
            .O(N__10728),
            .I(N__10725));
    Odrv4 I__2148 (
            .O(N__10725),
            .I(\d1.state_0_sqmuxaZ0Z_2 ));
    CascadeMux I__2147 (
            .O(N__10722),
            .I(\d1.state_0_sqmuxaZ0Z_2_cascade_ ));
    InMux I__2146 (
            .O(N__10719),
            .I(N__10716));
    LocalMux I__2145 (
            .O(N__10716),
            .I(state_0_sqmuxa));
    CascadeMux I__2144 (
            .O(N__10713),
            .I(state_0_sqmuxa_cascade_));
    InMux I__2143 (
            .O(N__10710),
            .I(N__10706));
    InMux I__2142 (
            .O(N__10709),
            .I(N__10703));
    LocalMux I__2141 (
            .O(N__10706),
            .I(N__10700));
    LocalMux I__2140 (
            .O(N__10703),
            .I(N__10697));
    Span4Mux_h I__2139 (
            .O(N__10700),
            .I(N__10694));
    Odrv4 I__2138 (
            .O(N__10697),
            .I(alarm_on_0_sqmuxa));
    Odrv4 I__2137 (
            .O(N__10694),
            .I(alarm_on_0_sqmuxa));
    InMux I__2136 (
            .O(N__10689),
            .I(N__10686));
    LocalMux I__2135 (
            .O(N__10686),
            .I(N__10683));
    Span4Mux_h I__2134 (
            .O(N__10683),
            .I(N__10679));
    InMux I__2133 (
            .O(N__10682),
            .I(N__10676));
    Span4Mux_h I__2132 (
            .O(N__10679),
            .I(N__10673));
    LocalMux I__2131 (
            .O(N__10676),
            .I(alarm_onZ0));
    Odrv4 I__2130 (
            .O(N__10673),
            .I(alarm_onZ0));
    InMux I__2129 (
            .O(N__10668),
            .I(N__10663));
    InMux I__2128 (
            .O(N__10667),
            .I(N__10660));
    InMux I__2127 (
            .O(N__10666),
            .I(N__10657));
    LocalMux I__2126 (
            .O(N__10663),
            .I(\d3.countZ0Z_16 ));
    LocalMux I__2125 (
            .O(N__10660),
            .I(\d3.countZ0Z_16 ));
    LocalMux I__2124 (
            .O(N__10657),
            .I(\d3.countZ0Z_16 ));
    InMux I__2123 (
            .O(N__10650),
            .I(N__10645));
    InMux I__2122 (
            .O(N__10649),
            .I(N__10642));
    InMux I__2121 (
            .O(N__10648),
            .I(N__10639));
    LocalMux I__2120 (
            .O(N__10645),
            .I(\d3.countZ0Z_15 ));
    LocalMux I__2119 (
            .O(N__10642),
            .I(\d3.countZ0Z_15 ));
    LocalMux I__2118 (
            .O(N__10639),
            .I(\d3.countZ0Z_15 ));
    InMux I__2117 (
            .O(N__10632),
            .I(N__10627));
    InMux I__2116 (
            .O(N__10631),
            .I(N__10624));
    InMux I__2115 (
            .O(N__10630),
            .I(N__10621));
    LocalMux I__2114 (
            .O(N__10627),
            .I(\d3.countZ0Z_14 ));
    LocalMux I__2113 (
            .O(N__10624),
            .I(\d3.countZ0Z_14 ));
    LocalMux I__2112 (
            .O(N__10621),
            .I(\d3.countZ0Z_14 ));
    InMux I__2111 (
            .O(N__10614),
            .I(N__10611));
    LocalMux I__2110 (
            .O(N__10611),
            .I(\d3.count_RNI4GDSZ0Z_16 ));
    InMux I__2109 (
            .O(N__10608),
            .I(N__10604));
    CascadeMux I__2108 (
            .O(N__10607),
            .I(N__10601));
    LocalMux I__2107 (
            .O(N__10604),
            .I(N__10596));
    InMux I__2106 (
            .O(N__10601),
            .I(N__10593));
    InMux I__2105 (
            .O(N__10600),
            .I(N__10590));
    InMux I__2104 (
            .O(N__10599),
            .I(N__10586));
    Span4Mux_v I__2103 (
            .O(N__10596),
            .I(N__10581));
    LocalMux I__2102 (
            .O(N__10593),
            .I(N__10581));
    LocalMux I__2101 (
            .O(N__10590),
            .I(N__10578));
    InMux I__2100 (
            .O(N__10589),
            .I(N__10575));
    LocalMux I__2099 (
            .O(N__10586),
            .I(N__10572));
    Span4Mux_h I__2098 (
            .O(N__10581),
            .I(N__10569));
    Odrv12 I__2097 (
            .O(N__10578),
            .I(ten_secsZ0Z_2));
    LocalMux I__2096 (
            .O(N__10575),
            .I(ten_secsZ0Z_2));
    Odrv4 I__2095 (
            .O(N__10572),
            .I(ten_secsZ0Z_2));
    Odrv4 I__2094 (
            .O(N__10569),
            .I(ten_secsZ0Z_2));
    IoInMux I__2093 (
            .O(N__10560),
            .I(N__10557));
    LocalMux I__2092 (
            .O(N__10557),
            .I(N__10554));
    Span4Mux_s3_h I__2091 (
            .O(N__10554),
            .I(N__10551));
    Span4Mux_h I__2090 (
            .O(N__10551),
            .I(N__10546));
    InMux I__2089 (
            .O(N__10550),
            .I(N__10541));
    InMux I__2088 (
            .O(N__10549),
            .I(N__10538));
    Span4Mux_h I__2087 (
            .O(N__10546),
            .I(N__10535));
    CascadeMux I__2086 (
            .O(N__10545),
            .I(N__10531));
    CascadeMux I__2085 (
            .O(N__10544),
            .I(N__10527));
    LocalMux I__2084 (
            .O(N__10541),
            .I(N__10524));
    LocalMux I__2083 (
            .O(N__10538),
            .I(N__10519));
    Span4Mux_h I__2082 (
            .O(N__10535),
            .I(N__10519));
    InMux I__2081 (
            .O(N__10534),
            .I(N__10516));
    InMux I__2080 (
            .O(N__10531),
            .I(N__10513));
    InMux I__2079 (
            .O(N__10530),
            .I(N__10510));
    InMux I__2078 (
            .O(N__10527),
            .I(N__10507));
    Odrv4 I__2077 (
            .O(N__10524),
            .I(un1_state_3));
    Odrv4 I__2076 (
            .O(N__10519),
            .I(un1_state_3));
    LocalMux I__2075 (
            .O(N__10516),
            .I(un1_state_3));
    LocalMux I__2074 (
            .O(N__10513),
            .I(un1_state_3));
    LocalMux I__2073 (
            .O(N__10510),
            .I(un1_state_3));
    LocalMux I__2072 (
            .O(N__10507),
            .I(un1_state_3));
    InMux I__2071 (
            .O(N__10494),
            .I(N__10491));
    LocalMux I__2070 (
            .O(N__10491),
            .I(N__10488));
    Span4Mux_h I__2069 (
            .O(N__10488),
            .I(N__10485));
    Odrv4 I__2068 (
            .O(N__10485),
            .I(\d1.g0_0Z0Z_2 ));
    InMux I__2067 (
            .O(N__10482),
            .I(N__10479));
    LocalMux I__2066 (
            .O(N__10479),
            .I(N__10475));
    InMux I__2065 (
            .O(N__10478),
            .I(N__10470));
    Span12Mux_v I__2064 (
            .O(N__10475),
            .I(N__10466));
    InMux I__2063 (
            .O(N__10474),
            .I(N__10461));
    InMux I__2062 (
            .O(N__10473),
            .I(N__10461));
    LocalMux I__2061 (
            .O(N__10470),
            .I(N__10458));
    InMux I__2060 (
            .O(N__10469),
            .I(N__10455));
    Odrv12 I__2059 (
            .O(N__10466),
            .I(secsZ0Z_2));
    LocalMux I__2058 (
            .O(N__10461),
            .I(secsZ0Z_2));
    Odrv4 I__2057 (
            .O(N__10458),
            .I(secsZ0Z_2));
    LocalMux I__2056 (
            .O(N__10455),
            .I(secsZ0Z_2));
    InMux I__2055 (
            .O(N__10446),
            .I(N__10443));
    LocalMux I__2054 (
            .O(N__10443),
            .I(N__10437));
    InMux I__2053 (
            .O(N__10442),
            .I(N__10432));
    InMux I__2052 (
            .O(N__10441),
            .I(N__10427));
    InMux I__2051 (
            .O(N__10440),
            .I(N__10427));
    Span12Mux_s9_h I__2050 (
            .O(N__10437),
            .I(N__10424));
    InMux I__2049 (
            .O(N__10436),
            .I(N__10421));
    InMux I__2048 (
            .O(N__10435),
            .I(N__10418));
    LocalMux I__2047 (
            .O(N__10432),
            .I(secsZ0Z_1));
    LocalMux I__2046 (
            .O(N__10427),
            .I(secsZ0Z_1));
    Odrv12 I__2045 (
            .O(N__10424),
            .I(secsZ0Z_1));
    LocalMux I__2044 (
            .O(N__10421),
            .I(secsZ0Z_1));
    LocalMux I__2043 (
            .O(N__10418),
            .I(secsZ0Z_1));
    InMux I__2042 (
            .O(N__10407),
            .I(N__10404));
    LocalMux I__2041 (
            .O(N__10404),
            .I(N__10401));
    Span4Mux_v I__2040 (
            .O(N__10401),
            .I(N__10395));
    CascadeMux I__2039 (
            .O(N__10400),
            .I(N__10392));
    CascadeMux I__2038 (
            .O(N__10399),
            .I(N__10389));
    InMux I__2037 (
            .O(N__10398),
            .I(N__10386));
    Sp12to4 I__2036 (
            .O(N__10395),
            .I(N__10383));
    InMux I__2035 (
            .O(N__10392),
            .I(N__10380));
    InMux I__2034 (
            .O(N__10389),
            .I(N__10377));
    LocalMux I__2033 (
            .O(N__10386),
            .I(secsZ0Z_3));
    Odrv12 I__2032 (
            .O(N__10383),
            .I(secsZ0Z_3));
    LocalMux I__2031 (
            .O(N__10380),
            .I(secsZ0Z_3));
    LocalMux I__2030 (
            .O(N__10377),
            .I(secsZ0Z_3));
    InMux I__2029 (
            .O(N__10368),
            .I(N__10365));
    LocalMux I__2028 (
            .O(N__10365),
            .I(N__10362));
    Span4Mux_v I__2027 (
            .O(N__10362),
            .I(N__10359));
    Span4Mux_h I__2026 (
            .O(N__10359),
            .I(N__10353));
    InMux I__2025 (
            .O(N__10358),
            .I(N__10343));
    InMux I__2024 (
            .O(N__10357),
            .I(N__10343));
    InMux I__2023 (
            .O(N__10356),
            .I(N__10343));
    Span4Mux_h I__2022 (
            .O(N__10353),
            .I(N__10340));
    InMux I__2021 (
            .O(N__10352),
            .I(N__10337));
    InMux I__2020 (
            .O(N__10351),
            .I(N__10332));
    InMux I__2019 (
            .O(N__10350),
            .I(N__10332));
    LocalMux I__2018 (
            .O(N__10343),
            .I(secsZ0Z_0));
    Odrv4 I__2017 (
            .O(N__10340),
            .I(secsZ0Z_0));
    LocalMux I__2016 (
            .O(N__10337),
            .I(secsZ0Z_0));
    LocalMux I__2015 (
            .O(N__10332),
            .I(secsZ0Z_0));
    InMux I__2014 (
            .O(N__10323),
            .I(N__10320));
    LocalMux I__2013 (
            .O(N__10320),
            .I(N__10316));
    InMux I__2012 (
            .O(N__10319),
            .I(N__10313));
    Odrv4 I__2011 (
            .O(N__10316),
            .I(decrement_time_0_secs9));
    LocalMux I__2010 (
            .O(N__10313),
            .I(decrement_time_0_secs9));
    InMux I__2009 (
            .O(N__10308),
            .I(\d2.un3_count_cry_10 ));
    InMux I__2008 (
            .O(N__10305),
            .I(\d2.un3_count_cry_11 ));
    InMux I__2007 (
            .O(N__10302),
            .I(\d2.un3_count_cry_12 ));
    InMux I__2006 (
            .O(N__10299),
            .I(\d2.un3_count_cry_13 ));
    InMux I__2005 (
            .O(N__10296),
            .I(\d2.un3_count_cry_14 ));
    InMux I__2004 (
            .O(N__10293),
            .I(\d2.un3_count_cry_15 ));
    SRMux I__2003 (
            .O(N__10290),
            .I(N__10281));
    SRMux I__2002 (
            .O(N__10289),
            .I(N__10281));
    SRMux I__2001 (
            .O(N__10288),
            .I(N__10281));
    GlobalMux I__2000 (
            .O(N__10281),
            .I(N__10278));
    gio2CtrlBuf I__1999 (
            .O(N__10278),
            .I(\d2.idle_i_g ));
    CEMux I__1998 (
            .O(N__10275),
            .I(N__10272));
    LocalMux I__1997 (
            .O(N__10272),
            .I(N__10269));
    Span4Mux_h I__1996 (
            .O(N__10269),
            .I(N__10266));
    Odrv4 I__1995 (
            .O(N__10266),
            .I(un1_state_0_sqmuxa_1_0_0));
    InMux I__1994 (
            .O(N__10263),
            .I(N__10260));
    LocalMux I__1993 (
            .O(N__10260),
            .I(N__10257));
    Odrv4 I__1992 (
            .O(N__10257),
            .I(\d1.state_1_sqmuxaZ0 ));
    InMux I__1991 (
            .O(N__10254),
            .I(N__10251));
    LocalMux I__1990 (
            .O(N__10251),
            .I(un1_state_0_sqmuxa_1_0));
    InMux I__1989 (
            .O(N__10248),
            .I(\d2.un3_count_cry_1 ));
    InMux I__1988 (
            .O(N__10245),
            .I(\d2.un3_count_cry_2 ));
    InMux I__1987 (
            .O(N__10242),
            .I(\d2.un3_count_cry_3 ));
    InMux I__1986 (
            .O(N__10239),
            .I(\d2.un3_count_cry_4 ));
    InMux I__1985 (
            .O(N__10236),
            .I(\d2.un3_count_cry_5 ));
    InMux I__1984 (
            .O(N__10233),
            .I(\d2.un3_count_cry_6 ));
    InMux I__1983 (
            .O(N__10230),
            .I(\d2.un3_count_cry_7 ));
    InMux I__1982 (
            .O(N__10227),
            .I(bfn_11_19_0_));
    InMux I__1981 (
            .O(N__10224),
            .I(\d2.un3_count_cry_9 ));
    InMux I__1980 (
            .O(N__10221),
            .I(N__10218));
    LocalMux I__1979 (
            .O(N__10218),
            .I(N__10214));
    InMux I__1978 (
            .O(N__10217),
            .I(N__10211));
    Odrv12 I__1977 (
            .O(N__10214),
            .I(\d1.trans_up_1_0 ));
    LocalMux I__1976 (
            .O(N__10211),
            .I(\d1.trans_up_1_0 ));
    CascadeMux I__1975 (
            .O(N__10206),
            .I(N__10203));
    InMux I__1974 (
            .O(N__10203),
            .I(N__10200));
    LocalMux I__1973 (
            .O(N__10200),
            .I(\d1.g2_i_a5_3 ));
    CascadeMux I__1972 (
            .O(N__10197),
            .I(\d1.g0_0_0Z0Z_1_cascade_ ));
    InMux I__1971 (
            .O(N__10194),
            .I(N__10191));
    LocalMux I__1970 (
            .O(N__10191),
            .I(\d1.g2Z0Z_10 ));
    CascadeMux I__1969 (
            .O(N__10188),
            .I(N__10184));
    InMux I__1968 (
            .O(N__10187),
            .I(N__10181));
    InMux I__1967 (
            .O(N__10184),
            .I(N__10178));
    LocalMux I__1966 (
            .O(N__10181),
            .I(N__10175));
    LocalMux I__1965 (
            .O(N__10178),
            .I(N__10172));
    Odrv4 I__1964 (
            .O(N__10175),
            .I(\d1.g0_2_0_a4Z0Z_2 ));
    Odrv4 I__1963 (
            .O(N__10172),
            .I(\d1.g0_2_0_a4Z0Z_2 ));
    InMux I__1962 (
            .O(N__10167),
            .I(N__10164));
    LocalMux I__1961 (
            .O(N__10164),
            .I(N__10158));
    InMux I__1960 (
            .O(N__10163),
            .I(N__10155));
    InMux I__1959 (
            .O(N__10162),
            .I(N__10150));
    InMux I__1958 (
            .O(N__10161),
            .I(N__10147));
    Span4Mux_v I__1957 (
            .O(N__10158),
            .I(N__10144));
    LocalMux I__1956 (
            .O(N__10155),
            .I(N__10141));
    InMux I__1955 (
            .O(N__10154),
            .I(N__10136));
    InMux I__1954 (
            .O(N__10153),
            .I(N__10136));
    LocalMux I__1953 (
            .O(N__10150),
            .I(s_dn));
    LocalMux I__1952 (
            .O(N__10147),
            .I(s_dn));
    Odrv4 I__1951 (
            .O(N__10144),
            .I(s_dn));
    Odrv4 I__1950 (
            .O(N__10141),
            .I(s_dn));
    LocalMux I__1949 (
            .O(N__10136),
            .I(s_dn));
    InMux I__1948 (
            .O(N__10125),
            .I(N__10121));
    InMux I__1947 (
            .O(N__10124),
            .I(N__10118));
    LocalMux I__1946 (
            .O(N__10121),
            .I(\d1.g0_2_0_o2_2 ));
    LocalMux I__1945 (
            .O(N__10118),
            .I(\d1.g0_2_0_o2_2 ));
    InMux I__1944 (
            .O(N__10113),
            .I(N__10110));
    LocalMux I__1943 (
            .O(N__10110),
            .I(N__10107));
    Odrv4 I__1942 (
            .O(N__10107),
            .I(\d1.g2_i_a5_0Z0Z_3 ));
    CascadeMux I__1941 (
            .O(N__10104),
            .I(\d1.g2_i_a5_0Z0Z_6_cascade_ ));
    InMux I__1940 (
            .O(N__10101),
            .I(N__10098));
    LocalMux I__1939 (
            .O(N__10098),
            .I(\d1.g2_i_a5Z0Z_2 ));
    InMux I__1938 (
            .O(N__10095),
            .I(N__10092));
    LocalMux I__1937 (
            .O(N__10092),
            .I(N__10089));
    Odrv4 I__1936 (
            .O(N__10089),
            .I(\d1.secs_0_sqmuxa_xZ0Z1 ));
    CascadeMux I__1935 (
            .O(N__10086),
            .I(N__10083));
    InMux I__1934 (
            .O(N__10083),
            .I(N__10080));
    LocalMux I__1933 (
            .O(N__10080),
            .I(N__10077));
    Span4Mux_h I__1932 (
            .O(N__10077),
            .I(N__10074));
    Span4Mux_h I__1931 (
            .O(N__10074),
            .I(N__10071));
    Odrv4 I__1930 (
            .O(N__10071),
            .I(mins_storedZ0Z_3));
    InMux I__1929 (
            .O(N__10068),
            .I(N__10065));
    LocalMux I__1928 (
            .O(N__10065),
            .I(\d1.N_5 ));
    InMux I__1927 (
            .O(N__10062),
            .I(N__10056));
    InMux I__1926 (
            .O(N__10061),
            .I(N__10053));
    InMux I__1925 (
            .O(N__10060),
            .I(N__10048));
    InMux I__1924 (
            .O(N__10059),
            .I(N__10048));
    LocalMux I__1923 (
            .O(N__10056),
            .I(\d1.un1_mins_1_sqmuxa_0 ));
    LocalMux I__1922 (
            .O(N__10053),
            .I(\d1.un1_mins_1_sqmuxa_0 ));
    LocalMux I__1921 (
            .O(N__10048),
            .I(\d1.un1_mins_1_sqmuxa_0 ));
    InMux I__1920 (
            .O(N__10041),
            .I(N__10038));
    LocalMux I__1919 (
            .O(N__10038),
            .I(N__10035));
    Odrv4 I__1918 (
            .O(N__10035),
            .I(\d1.g0_0_0_a4_2_1 ));
    CascadeMux I__1917 (
            .O(N__10032),
            .I(secs_RNO_0Z0Z_2_cascade_));
    InMux I__1916 (
            .O(N__10029),
            .I(N__10026));
    LocalMux I__1915 (
            .O(N__10026),
            .I(N__10020));
    InMux I__1914 (
            .O(N__10025),
            .I(N__10017));
    InMux I__1913 (
            .O(N__10024),
            .I(N__10014));
    InMux I__1912 (
            .O(N__10023),
            .I(N__10011));
    Odrv4 I__1911 (
            .O(N__10020),
            .I(secs_0_sqmuxa));
    LocalMux I__1910 (
            .O(N__10017),
            .I(secs_0_sqmuxa));
    LocalMux I__1909 (
            .O(N__10014),
            .I(secs_0_sqmuxa));
    LocalMux I__1908 (
            .O(N__10011),
            .I(secs_0_sqmuxa));
    CascadeMux I__1907 (
            .O(N__10002),
            .I(N__9996));
    CascadeMux I__1906 (
            .O(N__10001),
            .I(N__9993));
    InMux I__1905 (
            .O(N__10000),
            .I(N__9984));
    InMux I__1904 (
            .O(N__9999),
            .I(N__9984));
    InMux I__1903 (
            .O(N__9996),
            .I(N__9984));
    InMux I__1902 (
            .O(N__9993),
            .I(N__9984));
    LocalMux I__1901 (
            .O(N__9984),
            .I(un1_state_7_0));
    CascadeMux I__1900 (
            .O(N__9981),
            .I(un1_secs_c3_cascade_));
    InMux I__1899 (
            .O(N__9978),
            .I(N__9969));
    InMux I__1898 (
            .O(N__9977),
            .I(N__9969));
    InMux I__1897 (
            .O(N__9976),
            .I(N__9969));
    LocalMux I__1896 (
            .O(N__9969),
            .I(un1_alarm_on_0_sqmuxa_0_i));
    InMux I__1895 (
            .O(N__9966),
            .I(\d3.un3_count_cry_14 ));
    InMux I__1894 (
            .O(N__9963),
            .I(\d3.un3_count_cry_15 ));
    SRMux I__1893 (
            .O(N__9960),
            .I(N__9951));
    SRMux I__1892 (
            .O(N__9959),
            .I(N__9951));
    SRMux I__1891 (
            .O(N__9958),
            .I(N__9951));
    GlobalMux I__1890 (
            .O(N__9951),
            .I(N__9948));
    gio2CtrlBuf I__1889 (
            .O(N__9948),
            .I(\d3.idle_i_g ));
    InMux I__1888 (
            .O(N__9945),
            .I(N__9935));
    InMux I__1887 (
            .O(N__9944),
            .I(N__9920));
    InMux I__1886 (
            .O(N__9943),
            .I(N__9920));
    InMux I__1885 (
            .O(N__9942),
            .I(N__9920));
    InMux I__1884 (
            .O(N__9941),
            .I(N__9920));
    InMux I__1883 (
            .O(N__9940),
            .I(N__9920));
    InMux I__1882 (
            .O(N__9939),
            .I(N__9920));
    InMux I__1881 (
            .O(N__9938),
            .I(N__9920));
    LocalMux I__1880 (
            .O(N__9935),
            .I(N__9912));
    LocalMux I__1879 (
            .O(N__9920),
            .I(N__9908));
    InMux I__1878 (
            .O(N__9919),
            .I(N__9897));
    InMux I__1877 (
            .O(N__9918),
            .I(N__9897));
    InMux I__1876 (
            .O(N__9917),
            .I(N__9897));
    InMux I__1875 (
            .O(N__9916),
            .I(N__9897));
    InMux I__1874 (
            .O(N__9915),
            .I(N__9897));
    Span4Mux_h I__1873 (
            .O(N__9912),
            .I(N__9894));
    InMux I__1872 (
            .O(N__9911),
            .I(N__9891));
    Odrv4 I__1871 (
            .O(N__9908),
            .I(decrement_time_0_prescaler10_THRU_CO));
    LocalMux I__1870 (
            .O(N__9897),
            .I(decrement_time_0_prescaler10_THRU_CO));
    Odrv4 I__1869 (
            .O(N__9894),
            .I(decrement_time_0_prescaler10_THRU_CO));
    LocalMux I__1868 (
            .O(N__9891),
            .I(decrement_time_0_prescaler10_THRU_CO));
    CascadeMux I__1867 (
            .O(N__9882),
            .I(un1_state_7_0_cascade_));
    CascadeMux I__1866 (
            .O(N__9879),
            .I(un1_alarm_on_0_sqmuxa_0_i_cascade_));
    InMux I__1865 (
            .O(N__9876),
            .I(N__9873));
    LocalMux I__1864 (
            .O(N__9873),
            .I(N_120_1));
    InMux I__1863 (
            .O(N__9870),
            .I(N__9862));
    InMux I__1862 (
            .O(N__9869),
            .I(N__9859));
    InMux I__1861 (
            .O(N__9868),
            .I(N__9854));
    InMux I__1860 (
            .O(N__9867),
            .I(N__9854));
    InMux I__1859 (
            .O(N__9866),
            .I(N__9851));
    InMux I__1858 (
            .O(N__9865),
            .I(N__9848));
    LocalMux I__1857 (
            .O(N__9862),
            .I(s_cancel));
    LocalMux I__1856 (
            .O(N__9859),
            .I(s_cancel));
    LocalMux I__1855 (
            .O(N__9854),
            .I(s_cancel));
    LocalMux I__1854 (
            .O(N__9851),
            .I(s_cancel));
    LocalMux I__1853 (
            .O(N__9848),
            .I(s_cancel));
    CascadeMux I__1852 (
            .O(N__9837),
            .I(N__9833));
    InMux I__1851 (
            .O(N__9836),
            .I(N__9829));
    InMux I__1850 (
            .O(N__9833),
            .I(N__9826));
    InMux I__1849 (
            .O(N__9832),
            .I(N__9823));
    LocalMux I__1848 (
            .O(N__9829),
            .I(\d3.countZ0Z_13 ));
    LocalMux I__1847 (
            .O(N__9826),
            .I(\d3.countZ0Z_13 ));
    LocalMux I__1846 (
            .O(N__9823),
            .I(\d3.countZ0Z_13 ));
    InMux I__1845 (
            .O(N__9816),
            .I(N__9813));
    LocalMux I__1844 (
            .O(N__9813),
            .I(N__9809));
    InMux I__1843 (
            .O(N__9812),
            .I(N__9806));
    Odrv4 I__1842 (
            .O(N__9809),
            .I(d3_g0_1));
    LocalMux I__1841 (
            .O(N__9806),
            .I(d3_g0_1));
    InMux I__1840 (
            .O(N__9801),
            .I(N__9797));
    InMux I__1839 (
            .O(N__9800),
            .I(N__9794));
    LocalMux I__1838 (
            .O(N__9797),
            .I(\d3.countZ0Z_6 ));
    LocalMux I__1837 (
            .O(N__9794),
            .I(\d3.countZ0Z_6 ));
    InMux I__1836 (
            .O(N__9789),
            .I(\d3.un3_count_cry_5 ));
    InMux I__1835 (
            .O(N__9786),
            .I(N__9782));
    InMux I__1834 (
            .O(N__9785),
            .I(N__9779));
    LocalMux I__1833 (
            .O(N__9782),
            .I(\d3.countZ0Z_7 ));
    LocalMux I__1832 (
            .O(N__9779),
            .I(\d3.countZ0Z_7 ));
    InMux I__1831 (
            .O(N__9774),
            .I(\d3.un3_count_cry_6 ));
    InMux I__1830 (
            .O(N__9771),
            .I(N__9767));
    InMux I__1829 (
            .O(N__9770),
            .I(N__9764));
    LocalMux I__1828 (
            .O(N__9767),
            .I(\d3.countZ0Z_8 ));
    LocalMux I__1827 (
            .O(N__9764),
            .I(\d3.countZ0Z_8 ));
    InMux I__1826 (
            .O(N__9759),
            .I(\d3.un3_count_cry_7 ));
    CascadeMux I__1825 (
            .O(N__9756),
            .I(N__9752));
    InMux I__1824 (
            .O(N__9755),
            .I(N__9749));
    InMux I__1823 (
            .O(N__9752),
            .I(N__9746));
    LocalMux I__1822 (
            .O(N__9749),
            .I(\d3.countZ0Z_9 ));
    LocalMux I__1821 (
            .O(N__9746),
            .I(\d3.countZ0Z_9 ));
    InMux I__1820 (
            .O(N__9741),
            .I(bfn_11_14_0_));
    InMux I__1819 (
            .O(N__9738),
            .I(N__9734));
    InMux I__1818 (
            .O(N__9737),
            .I(N__9731));
    LocalMux I__1817 (
            .O(N__9734),
            .I(N__9728));
    LocalMux I__1816 (
            .O(N__9731),
            .I(\d3.countZ0Z_10 ));
    Odrv4 I__1815 (
            .O(N__9728),
            .I(\d3.countZ0Z_10 ));
    InMux I__1814 (
            .O(N__9723),
            .I(\d3.un3_count_cry_9 ));
    CascadeMux I__1813 (
            .O(N__9720),
            .I(N__9717));
    InMux I__1812 (
            .O(N__9717),
            .I(N__9713));
    InMux I__1811 (
            .O(N__9716),
            .I(N__9710));
    LocalMux I__1810 (
            .O(N__9713),
            .I(N__9707));
    LocalMux I__1809 (
            .O(N__9710),
            .I(\d3.countZ0Z_11 ));
    Odrv4 I__1808 (
            .O(N__9707),
            .I(\d3.countZ0Z_11 ));
    InMux I__1807 (
            .O(N__9702),
            .I(\d3.un3_count_cry_10 ));
    CascadeMux I__1806 (
            .O(N__9699),
            .I(N__9696));
    InMux I__1805 (
            .O(N__9696),
            .I(N__9692));
    InMux I__1804 (
            .O(N__9695),
            .I(N__9689));
    LocalMux I__1803 (
            .O(N__9692),
            .I(N__9686));
    LocalMux I__1802 (
            .O(N__9689),
            .I(\d3.countZ0Z_12 ));
    Odrv12 I__1801 (
            .O(N__9686),
            .I(\d3.countZ0Z_12 ));
    InMux I__1800 (
            .O(N__9681),
            .I(\d3.un3_count_cry_11 ));
    InMux I__1799 (
            .O(N__9678),
            .I(\d3.un3_count_cry_12 ));
    InMux I__1798 (
            .O(N__9675),
            .I(\d3.un3_count_cry_13 ));
    CascadeMux I__1797 (
            .O(N__9672),
            .I(N__9668));
    InMux I__1796 (
            .O(N__9671),
            .I(N__9665));
    InMux I__1795 (
            .O(N__9668),
            .I(N__9662));
    LocalMux I__1794 (
            .O(N__9665),
            .I(\d4.countZ0Z_14 ));
    LocalMux I__1793 (
            .O(N__9662),
            .I(\d4.countZ0Z_14 ));
    InMux I__1792 (
            .O(N__9657),
            .I(\d4.un3_count_cry_13 ));
    InMux I__1791 (
            .O(N__9654),
            .I(N__9650));
    InMux I__1790 (
            .O(N__9653),
            .I(N__9647));
    LocalMux I__1789 (
            .O(N__9650),
            .I(\d4.countZ0Z_15 ));
    LocalMux I__1788 (
            .O(N__9647),
            .I(\d4.countZ0Z_15 ));
    InMux I__1787 (
            .O(N__9642),
            .I(\d4.un3_count_cry_14 ));
    InMux I__1786 (
            .O(N__9639),
            .I(\d4.un3_count_cry_15 ));
    CascadeMux I__1785 (
            .O(N__9636),
            .I(N__9632));
    InMux I__1784 (
            .O(N__9635),
            .I(N__9629));
    InMux I__1783 (
            .O(N__9632),
            .I(N__9626));
    LocalMux I__1782 (
            .O(N__9629),
            .I(\d4.countZ0Z_16 ));
    LocalMux I__1781 (
            .O(N__9626),
            .I(\d4.countZ0Z_16 ));
    SRMux I__1780 (
            .O(N__9621),
            .I(N__9612));
    SRMux I__1779 (
            .O(N__9620),
            .I(N__9612));
    SRMux I__1778 (
            .O(N__9619),
            .I(N__9612));
    GlobalMux I__1777 (
            .O(N__9612),
            .I(N__9609));
    gio2CtrlBuf I__1776 (
            .O(N__9609),
            .I(\d4.idle_i_g ));
    InMux I__1775 (
            .O(N__9606),
            .I(N__9600));
    InMux I__1774 (
            .O(N__9605),
            .I(N__9593));
    InMux I__1773 (
            .O(N__9604),
            .I(N__9593));
    InMux I__1772 (
            .O(N__9603),
            .I(N__9593));
    LocalMux I__1771 (
            .O(N__9600),
            .I(\d3.countZ0Z_0 ));
    LocalMux I__1770 (
            .O(N__9593),
            .I(\d3.countZ0Z_0 ));
    CascadeMux I__1769 (
            .O(N__9588),
            .I(N__9584));
    CascadeMux I__1768 (
            .O(N__9587),
            .I(N__9581));
    InMux I__1767 (
            .O(N__9584),
            .I(N__9577));
    InMux I__1766 (
            .O(N__9581),
            .I(N__9572));
    InMux I__1765 (
            .O(N__9580),
            .I(N__9572));
    LocalMux I__1764 (
            .O(N__9577),
            .I(\d3.countZ0Z_1 ));
    LocalMux I__1763 (
            .O(N__9572),
            .I(\d3.countZ0Z_1 ));
    InMux I__1762 (
            .O(N__9567),
            .I(N__9563));
    InMux I__1761 (
            .O(N__9566),
            .I(N__9560));
    LocalMux I__1760 (
            .O(N__9563),
            .I(\d3.countZ0Z_2 ));
    LocalMux I__1759 (
            .O(N__9560),
            .I(\d3.countZ0Z_2 ));
    InMux I__1758 (
            .O(N__9555),
            .I(\d3.un3_count_cry_1 ));
    InMux I__1757 (
            .O(N__9552),
            .I(N__9548));
    InMux I__1756 (
            .O(N__9551),
            .I(N__9545));
    LocalMux I__1755 (
            .O(N__9548),
            .I(\d3.countZ0Z_3 ));
    LocalMux I__1754 (
            .O(N__9545),
            .I(\d3.countZ0Z_3 ));
    InMux I__1753 (
            .O(N__9540),
            .I(\d3.un3_count_cry_2 ));
    InMux I__1752 (
            .O(N__9537),
            .I(N__9533));
    InMux I__1751 (
            .O(N__9536),
            .I(N__9530));
    LocalMux I__1750 (
            .O(N__9533),
            .I(\d3.countZ0Z_4 ));
    LocalMux I__1749 (
            .O(N__9530),
            .I(\d3.countZ0Z_4 ));
    InMux I__1748 (
            .O(N__9525),
            .I(\d3.un3_count_cry_3 ));
    CascadeMux I__1747 (
            .O(N__9522),
            .I(N__9518));
    InMux I__1746 (
            .O(N__9521),
            .I(N__9515));
    InMux I__1745 (
            .O(N__9518),
            .I(N__9512));
    LocalMux I__1744 (
            .O(N__9515),
            .I(\d3.countZ0Z_5 ));
    LocalMux I__1743 (
            .O(N__9512),
            .I(\d3.countZ0Z_5 ));
    InMux I__1742 (
            .O(N__9507),
            .I(\d3.un3_count_cry_4 ));
    InMux I__1741 (
            .O(N__9504),
            .I(\d4.un3_count_cry_4 ));
    CascadeMux I__1740 (
            .O(N__9501),
            .I(N__9497));
    InMux I__1739 (
            .O(N__9500),
            .I(N__9494));
    InMux I__1738 (
            .O(N__9497),
            .I(N__9491));
    LocalMux I__1737 (
            .O(N__9494),
            .I(\d4.countZ0Z_6 ));
    LocalMux I__1736 (
            .O(N__9491),
            .I(\d4.countZ0Z_6 ));
    InMux I__1735 (
            .O(N__9486),
            .I(\d4.un3_count_cry_5 ));
    InMux I__1734 (
            .O(N__9483),
            .I(N__9479));
    InMux I__1733 (
            .O(N__9482),
            .I(N__9476));
    LocalMux I__1732 (
            .O(N__9479),
            .I(\d4.countZ0Z_7 ));
    LocalMux I__1731 (
            .O(N__9476),
            .I(\d4.countZ0Z_7 ));
    InMux I__1730 (
            .O(N__9471),
            .I(\d4.un3_count_cry_6 ));
    InMux I__1729 (
            .O(N__9468),
            .I(N__9464));
    InMux I__1728 (
            .O(N__9467),
            .I(N__9461));
    LocalMux I__1727 (
            .O(N__9464),
            .I(\d4.countZ0Z_8 ));
    LocalMux I__1726 (
            .O(N__9461),
            .I(\d4.countZ0Z_8 ));
    InMux I__1725 (
            .O(N__9456),
            .I(\d4.un3_count_cry_7 ));
    InMux I__1724 (
            .O(N__9453),
            .I(N__9449));
    InMux I__1723 (
            .O(N__9452),
            .I(N__9446));
    LocalMux I__1722 (
            .O(N__9449),
            .I(\d4.countZ0Z_9 ));
    LocalMux I__1721 (
            .O(N__9446),
            .I(\d4.countZ0Z_9 ));
    InMux I__1720 (
            .O(N__9441),
            .I(bfn_11_12_0_));
    CascadeMux I__1719 (
            .O(N__9438),
            .I(N__9434));
    InMux I__1718 (
            .O(N__9437),
            .I(N__9431));
    InMux I__1717 (
            .O(N__9434),
            .I(N__9428));
    LocalMux I__1716 (
            .O(N__9431),
            .I(\d4.countZ0Z_10 ));
    LocalMux I__1715 (
            .O(N__9428),
            .I(\d4.countZ0Z_10 ));
    InMux I__1714 (
            .O(N__9423),
            .I(\d4.un3_count_cry_9 ));
    InMux I__1713 (
            .O(N__9420),
            .I(N__9416));
    InMux I__1712 (
            .O(N__9419),
            .I(N__9413));
    LocalMux I__1711 (
            .O(N__9416),
            .I(\d4.countZ0Z_11 ));
    LocalMux I__1710 (
            .O(N__9413),
            .I(\d4.countZ0Z_11 ));
    InMux I__1709 (
            .O(N__9408),
            .I(\d4.un3_count_cry_10 ));
    CascadeMux I__1708 (
            .O(N__9405),
            .I(N__9401));
    InMux I__1707 (
            .O(N__9404),
            .I(N__9398));
    InMux I__1706 (
            .O(N__9401),
            .I(N__9395));
    LocalMux I__1705 (
            .O(N__9398),
            .I(\d4.countZ0Z_12 ));
    LocalMux I__1704 (
            .O(N__9395),
            .I(\d4.countZ0Z_12 ));
    InMux I__1703 (
            .O(N__9390),
            .I(\d4.un3_count_cry_11 ));
    InMux I__1702 (
            .O(N__9387),
            .I(N__9383));
    InMux I__1701 (
            .O(N__9386),
            .I(N__9380));
    LocalMux I__1700 (
            .O(N__9383),
            .I(\d4.countZ0Z_13 ));
    LocalMux I__1699 (
            .O(N__9380),
            .I(\d4.countZ0Z_13 ));
    InMux I__1698 (
            .O(N__9375),
            .I(\d4.un3_count_cry_12 ));
    CascadeMux I__1697 (
            .O(N__9372),
            .I(\d1.g2Z0Z_7_cascade_ ));
    CascadeMux I__1696 (
            .O(N__9369),
            .I(\d1.g0_1_0_a4Z0Z_7_cascade_ ));
    InMux I__1695 (
            .O(N__9366),
            .I(N__9363));
    LocalMux I__1694 (
            .O(N__9363),
            .I(N__9357));
    InMux I__1693 (
            .O(N__9362),
            .I(N__9352));
    InMux I__1692 (
            .O(N__9361),
            .I(N__9352));
    InMux I__1691 (
            .O(N__9360),
            .I(N__9349));
    Span4Mux_v I__1690 (
            .O(N__9357),
            .I(N__9346));
    LocalMux I__1689 (
            .O(N__9352),
            .I(\d4.countZ0Z_0 ));
    LocalMux I__1688 (
            .O(N__9349),
            .I(\d4.countZ0Z_0 ));
    Odrv4 I__1687 (
            .O(N__9346),
            .I(\d4.countZ0Z_0 ));
    CascadeMux I__1686 (
            .O(N__9339),
            .I(N__9334));
    InMux I__1685 (
            .O(N__9338),
            .I(N__9331));
    InMux I__1684 (
            .O(N__9337),
            .I(N__9328));
    InMux I__1683 (
            .O(N__9334),
            .I(N__9325));
    LocalMux I__1682 (
            .O(N__9331),
            .I(N__9322));
    LocalMux I__1681 (
            .O(N__9328),
            .I(\d4.countZ0Z_1 ));
    LocalMux I__1680 (
            .O(N__9325),
            .I(\d4.countZ0Z_1 ));
    Odrv4 I__1679 (
            .O(N__9322),
            .I(\d4.countZ0Z_1 ));
    InMux I__1678 (
            .O(N__9315),
            .I(N__9311));
    InMux I__1677 (
            .O(N__9314),
            .I(N__9308));
    LocalMux I__1676 (
            .O(N__9311),
            .I(\d4.countZ0Z_2 ));
    LocalMux I__1675 (
            .O(N__9308),
            .I(\d4.countZ0Z_2 ));
    InMux I__1674 (
            .O(N__9303),
            .I(\d4.un3_count_cry_1 ));
    InMux I__1673 (
            .O(N__9300),
            .I(N__9296));
    InMux I__1672 (
            .O(N__9299),
            .I(N__9293));
    LocalMux I__1671 (
            .O(N__9296),
            .I(\d4.countZ0Z_3 ));
    LocalMux I__1670 (
            .O(N__9293),
            .I(\d4.countZ0Z_3 ));
    InMux I__1669 (
            .O(N__9288),
            .I(\d4.un3_count_cry_2 ));
    InMux I__1668 (
            .O(N__9285),
            .I(N__9281));
    InMux I__1667 (
            .O(N__9284),
            .I(N__9278));
    LocalMux I__1666 (
            .O(N__9281),
            .I(\d4.countZ0Z_4 ));
    LocalMux I__1665 (
            .O(N__9278),
            .I(\d4.countZ0Z_4 ));
    InMux I__1664 (
            .O(N__9273),
            .I(\d4.un3_count_cry_3 ));
    InMux I__1663 (
            .O(N__9270),
            .I(N__9266));
    InMux I__1662 (
            .O(N__9269),
            .I(N__9263));
    LocalMux I__1661 (
            .O(N__9266),
            .I(\d4.countZ0Z_5 ));
    LocalMux I__1660 (
            .O(N__9263),
            .I(\d4.countZ0Z_5 ));
    InMux I__1659 (
            .O(N__9258),
            .I(N__9255));
    LocalMux I__1658 (
            .O(N__9255),
            .I(N__9252));
    Odrv4 I__1657 (
            .O(N__9252),
            .I(\d1.g2_8_1 ));
    CascadeMux I__1656 (
            .O(N__9249),
            .I(\d2.g0_0_10_cascade_ ));
    InMux I__1655 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__1654 (
            .O(N__9243),
            .I(\d2.g0_0_12 ));
    CascadeMux I__1653 (
            .O(N__9240),
            .I(\d2.g0_0_14_cascade_ ));
    InMux I__1652 (
            .O(N__9237),
            .I(N__9234));
    LocalMux I__1651 (
            .O(N__9234),
            .I(N__9231));
    Odrv4 I__1650 (
            .O(N__9231),
            .I(\d1.g2_8_0 ));
    InMux I__1649 (
            .O(N__9228),
            .I(N__9225));
    LocalMux I__1648 (
            .O(N__9225),
            .I(\d2.g0_0_11 ));
    CascadeMux I__1647 (
            .O(N__9222),
            .I(N__9219));
    InMux I__1646 (
            .O(N__9219),
            .I(N__9216));
    LocalMux I__1645 (
            .O(N__9216),
            .I(\d2.trans_up_1_14_2 ));
    InMux I__1644 (
            .O(N__9213),
            .I(N__9210));
    LocalMux I__1643 (
            .O(N__9210),
            .I(\d1.g1_7 ));
    CascadeMux I__1642 (
            .O(N__9207),
            .I(N__9204));
    InMux I__1641 (
            .O(N__9204),
            .I(N__9201));
    LocalMux I__1640 (
            .O(N__9201),
            .I(\d1.g1_8 ));
    InMux I__1639 (
            .O(N__9198),
            .I(N__9195));
    LocalMux I__1638 (
            .O(N__9195),
            .I(\d1.g1_14 ));
    InMux I__1637 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__1636 (
            .O(N__9189),
            .I(N__9186));
    Span4Mux_h I__1635 (
            .O(N__9186),
            .I(N__9183));
    Odrv4 I__1634 (
            .O(N__9183),
            .I(\d1.g0_1_a5_0_10 ));
    InMux I__1633 (
            .O(N__9180),
            .I(N__9177));
    LocalMux I__1632 (
            .O(N__9177),
            .I(N__9174));
    Odrv4 I__1631 (
            .O(N__9174),
            .I(\d1.g0_1_a5_0_15 ));
    InMux I__1630 (
            .O(N__9171),
            .I(N__9168));
    LocalMux I__1629 (
            .O(N__9168),
            .I(N__9164));
    InMux I__1628 (
            .O(N__9167),
            .I(N__9161));
    Span4Mux_h I__1627 (
            .O(N__9164),
            .I(N__9158));
    LocalMux I__1626 (
            .O(N__9161),
            .I(\d1.trans_up_1_10 ));
    Odrv4 I__1625 (
            .O(N__9158),
            .I(\d1.trans_up_1_10 ));
    CascadeMux I__1624 (
            .O(N__9153),
            .I(N__9149));
    InMux I__1623 (
            .O(N__9152),
            .I(N__9146));
    InMux I__1622 (
            .O(N__9149),
            .I(N__9143));
    LocalMux I__1621 (
            .O(N__9146),
            .I(N__9140));
    LocalMux I__1620 (
            .O(N__9143),
            .I(N__9137));
    Span4Mux_v I__1619 (
            .O(N__9140),
            .I(N__9132));
    Span4Mux_h I__1618 (
            .O(N__9137),
            .I(N__9132));
    Span4Mux_h I__1617 (
            .O(N__9132),
            .I(N__9129));
    Odrv4 I__1616 (
            .O(N__9129),
            .I(\d1.trans_up_1_11 ));
    InMux I__1615 (
            .O(N__9126),
            .I(N__9123));
    LocalMux I__1614 (
            .O(N__9123),
            .I(N__9120));
    Span4Mux_v I__1613 (
            .O(N__9120),
            .I(N__9116));
    InMux I__1612 (
            .O(N__9119),
            .I(N__9113));
    Odrv4 I__1611 (
            .O(N__9116),
            .I(\d1.trans_up_1_13 ));
    LocalMux I__1610 (
            .O(N__9113),
            .I(\d1.trans_up_1_13 ));
    CascadeMux I__1609 (
            .O(N__9108),
            .I(\d1.trans_up_1_0_cascade_ ));
    CascadeMux I__1608 (
            .O(N__9105),
            .I(\d1.g0_2_0_o2_2_cascade_ ));
    InMux I__1607 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__1606 (
            .O(N__9099),
            .I(N__9096));
    Span4Mux_h I__1605 (
            .O(N__9096),
            .I(N__9093));
    Odrv4 I__1604 (
            .O(N__9093),
            .I(mins_storedZ0Z_0));
    InMux I__1603 (
            .O(N__9090),
            .I(N__9087));
    LocalMux I__1602 (
            .O(N__9087),
            .I(\d1.g0_0_0 ));
    CascadeMux I__1601 (
            .O(N__9084),
            .I(\d1.N_19_i_cascade_ ));
    CascadeMux I__1600 (
            .O(N__9081),
            .I(N__9077));
    InMux I__1599 (
            .O(N__9080),
            .I(N__9073));
    InMux I__1598 (
            .O(N__9077),
            .I(N__9070));
    CascadeMux I__1597 (
            .O(N__9076),
            .I(N__9067));
    LocalMux I__1596 (
            .O(N__9073),
            .I(N__9060));
    LocalMux I__1595 (
            .O(N__9070),
            .I(N__9060));
    InMux I__1594 (
            .O(N__9067),
            .I(N__9057));
    CascadeMux I__1593 (
            .O(N__9066),
            .I(N__9053));
    InMux I__1592 (
            .O(N__9065),
            .I(N__9049));
    Span4Mux_h I__1591 (
            .O(N__9060),
            .I(N__9043));
    LocalMux I__1590 (
            .O(N__9057),
            .I(N__9043));
    InMux I__1589 (
            .O(N__9056),
            .I(N__9038));
    InMux I__1588 (
            .O(N__9053),
            .I(N__9038));
    InMux I__1587 (
            .O(N__9052),
            .I(N__9035));
    LocalMux I__1586 (
            .O(N__9049),
            .I(N__9032));
    InMux I__1585 (
            .O(N__9048),
            .I(N__9029));
    Span4Mux_h I__1584 (
            .O(N__9043),
            .I(N__9026));
    LocalMux I__1583 (
            .O(N__9038),
            .I(N__9023));
    LocalMux I__1582 (
            .O(N__9035),
            .I(\d1.stateZ0Z_0 ));
    Odrv12 I__1581 (
            .O(N__9032),
            .I(\d1.stateZ0Z_0 ));
    LocalMux I__1580 (
            .O(N__9029),
            .I(\d1.stateZ0Z_0 ));
    Odrv4 I__1579 (
            .O(N__9026),
            .I(\d1.stateZ0Z_0 ));
    Odrv4 I__1578 (
            .O(N__9023),
            .I(\d1.stateZ0Z_0 ));
    CascadeMux I__1577 (
            .O(N__9012),
            .I(N__9009));
    InMux I__1576 (
            .O(N__9009),
            .I(N__9006));
    LocalMux I__1575 (
            .O(N__9006),
            .I(N__9003));
    Odrv12 I__1574 (
            .O(N__9003),
            .I(\d1.ten_secs_1_sqmuxa_0 ));
    InMux I__1573 (
            .O(N__9000),
            .I(N__8997));
    LocalMux I__1572 (
            .O(N__8997),
            .I(\d1.g2_0Z0Z_4 ));
    InMux I__1571 (
            .O(N__8994),
            .I(N__8991));
    LocalMux I__1570 (
            .O(N__8991),
            .I(N__8988));
    Odrv12 I__1569 (
            .O(N__8988),
            .I(\d1.g2_0Z0Z_3 ));
    CascadeMux I__1568 (
            .O(N__8985),
            .I(ten_secs_1_sqmuxa_cascade_));
    InMux I__1567 (
            .O(N__8982),
            .I(N__8979));
    LocalMux I__1566 (
            .O(N__8979),
            .I(N__8976));
    Odrv12 I__1565 (
            .O(N__8976),
            .I(\d1.g1_0 ));
    CascadeMux I__1564 (
            .O(N__8973),
            .I(\d1.g0_0_0_0_0_cascade_ ));
    InMux I__1563 (
            .O(N__8970),
            .I(N__8967));
    LocalMux I__1562 (
            .O(N__8967),
            .I(mins_storedZ0Z_1));
    CascadeMux I__1561 (
            .O(N__8964),
            .I(\d1.un1_mins_4_0_1_cascade_ ));
    InMux I__1560 (
            .O(N__8961),
            .I(N__8957));
    InMux I__1559 (
            .O(N__8960),
            .I(N__8953));
    LocalMux I__1558 (
            .O(N__8957),
            .I(N__8950));
    InMux I__1557 (
            .O(N__8956),
            .I(N__8947));
    LocalMux I__1556 (
            .O(N__8953),
            .I(N__8944));
    Span4Mux_h I__1555 (
            .O(N__8950),
            .I(N__8941));
    LocalMux I__1554 (
            .O(N__8947),
            .I(\d1.countZ0Z_9 ));
    Odrv12 I__1553 (
            .O(N__8944),
            .I(\d1.countZ0Z_9 ));
    Odrv4 I__1552 (
            .O(N__8941),
            .I(\d1.countZ0Z_9 ));
    InMux I__1551 (
            .O(N__8934),
            .I(N__8930));
    InMux I__1550 (
            .O(N__8933),
            .I(N__8926));
    LocalMux I__1549 (
            .O(N__8930),
            .I(N__8923));
    InMux I__1548 (
            .O(N__8929),
            .I(N__8920));
    LocalMux I__1547 (
            .O(N__8926),
            .I(N__8917));
    Span4Mux_h I__1546 (
            .O(N__8923),
            .I(N__8914));
    LocalMux I__1545 (
            .O(N__8920),
            .I(\d1.countZ0Z_8 ));
    Odrv12 I__1544 (
            .O(N__8917),
            .I(\d1.countZ0Z_8 ));
    Odrv4 I__1543 (
            .O(N__8914),
            .I(\d1.countZ0Z_8 ));
    CascadeMux I__1542 (
            .O(N__8907),
            .I(N__8904));
    InMux I__1541 (
            .O(N__8904),
            .I(N__8900));
    InMux I__1540 (
            .O(N__8903),
            .I(N__8896));
    LocalMux I__1539 (
            .O(N__8900),
            .I(N__8893));
    InMux I__1538 (
            .O(N__8899),
            .I(N__8890));
    LocalMux I__1537 (
            .O(N__8896),
            .I(N__8887));
    Span4Mux_h I__1536 (
            .O(N__8893),
            .I(N__8884));
    LocalMux I__1535 (
            .O(N__8890),
            .I(\d1.countZ0Z_10 ));
    Odrv12 I__1534 (
            .O(N__8887),
            .I(\d1.countZ0Z_10 ));
    Odrv4 I__1533 (
            .O(N__8884),
            .I(\d1.countZ0Z_10 ));
    InMux I__1532 (
            .O(N__8877),
            .I(N__8872));
    InMux I__1531 (
            .O(N__8876),
            .I(N__8869));
    InMux I__1530 (
            .O(N__8875),
            .I(N__8866));
    LocalMux I__1529 (
            .O(N__8872),
            .I(N__8863));
    LocalMux I__1528 (
            .O(N__8869),
            .I(N__8858));
    LocalMux I__1527 (
            .O(N__8866),
            .I(N__8858));
    Span4Mux_h I__1526 (
            .O(N__8863),
            .I(N__8855));
    Odrv4 I__1525 (
            .O(N__8858),
            .I(\d1.countZ0Z_7 ));
    Odrv4 I__1524 (
            .O(N__8855),
            .I(\d1.countZ0Z_7 ));
    InMux I__1523 (
            .O(N__8850),
            .I(N__8846));
    InMux I__1522 (
            .O(N__8849),
            .I(N__8843));
    LocalMux I__1521 (
            .O(N__8846),
            .I(\d1.trans_up_1_9 ));
    LocalMux I__1520 (
            .O(N__8843),
            .I(\d1.trans_up_1_9 ));
    InMux I__1519 (
            .O(N__8838),
            .I(N__8835));
    LocalMux I__1518 (
            .O(N__8835),
            .I(\d1.g2Z0Z_11 ));
    CascadeMux I__1517 (
            .O(N__8832),
            .I(\d1.un1_mins_1_sqmuxa_0_cascade_ ));
    CascadeMux I__1516 (
            .O(N__8829),
            .I(\d1.un1_mins_3_sqmuxa_0_0_cascade_ ));
    InMux I__1515 (
            .O(N__8826),
            .I(N__8823));
    LocalMux I__1514 (
            .O(N__8823),
            .I(\d1.N_4 ));
    InMux I__1513 (
            .O(N__8820),
            .I(N__8817));
    LocalMux I__1512 (
            .O(N__8817),
            .I(N__8814));
    Odrv4 I__1511 (
            .O(N__8814),
            .I(mins_storedZ0Z_2));
    CascadeMux I__1510 (
            .O(N__8811),
            .I(\d1.g1_cascade_ ));
    CascadeMux I__1509 (
            .O(N__8808),
            .I(d4_trans_up_1_cascade_));
    CascadeMux I__1508 (
            .O(N__8805),
            .I(ten_secs_r_1_1_cascade_));
    CascadeMux I__1507 (
            .O(N__8802),
            .I(\d3.trans_up_1_14_2_cascade_ ));
    CascadeMux I__1506 (
            .O(N__8799),
            .I(s_cancel_cascade_));
    InMux I__1505 (
            .O(N__8796),
            .I(N__8789));
    InMux I__1504 (
            .O(N__8795),
            .I(N__8786));
    InMux I__1503 (
            .O(N__8794),
            .I(N__8779));
    InMux I__1502 (
            .O(N__8793),
            .I(N__8779));
    InMux I__1501 (
            .O(N__8792),
            .I(N__8779));
    LocalMux I__1500 (
            .O(N__8789),
            .I(N__8776));
    LocalMux I__1499 (
            .O(N__8786),
            .I(N__8773));
    LocalMux I__1498 (
            .O(N__8779),
            .I(N__8770));
    Odrv4 I__1497 (
            .O(N__8776),
            .I(d4_state));
    Odrv12 I__1496 (
            .O(N__8773),
            .I(d4_state));
    Odrv4 I__1495 (
            .O(N__8770),
            .I(d4_state));
    InMux I__1494 (
            .O(N__8763),
            .I(N__8759));
    InMux I__1493 (
            .O(N__8762),
            .I(N__8756));
    LocalMux I__1492 (
            .O(N__8759),
            .I(d4_trans_up_1));
    LocalMux I__1491 (
            .O(N__8756),
            .I(d4_trans_up_1));
    CascadeMux I__1490 (
            .O(N__8751),
            .I(secs_0_sqmuxa_cascade_));
    InMux I__1489 (
            .O(N__8748),
            .I(N__8744));
    InMux I__1488 (
            .O(N__8747),
            .I(N__8740));
    LocalMux I__1487 (
            .O(N__8744),
            .I(N__8737));
    InMux I__1486 (
            .O(N__8743),
            .I(N__8734));
    LocalMux I__1485 (
            .O(N__8740),
            .I(un1_state_9_0));
    Odrv4 I__1484 (
            .O(N__8737),
            .I(un1_state_9_0));
    LocalMux I__1483 (
            .O(N__8734),
            .I(un1_state_9_0));
    InMux I__1482 (
            .O(N__8727),
            .I(N__8724));
    LocalMux I__1481 (
            .O(N__8724),
            .I(\d3.trans_up_1_15_8 ));
    InMux I__1480 (
            .O(N__8721),
            .I(N__8717));
    InMux I__1479 (
            .O(N__8720),
            .I(N__8714));
    LocalMux I__1478 (
            .O(N__8717),
            .I(N__8709));
    LocalMux I__1477 (
            .O(N__8714),
            .I(N__8709));
    Odrv12 I__1476 (
            .O(N__8709),
            .I(\d4.syncZ0Z_1 ));
    InMux I__1475 (
            .O(N__8706),
            .I(N__8703));
    LocalMux I__1474 (
            .O(N__8703),
            .I(\d3.trans_up_1_15_7 ));
    InMux I__1473 (
            .O(N__8700),
            .I(N__8697));
    LocalMux I__1472 (
            .O(N__8697),
            .I(N__8694));
    Odrv4 I__1471 (
            .O(N__8694),
            .I(\d4.trans_up_1_9 ));
    InMux I__1470 (
            .O(N__8691),
            .I(N__8688));
    LocalMux I__1469 (
            .O(N__8688),
            .I(\d4.trans_up_1_12 ));
    InMux I__1468 (
            .O(N__8685),
            .I(N__8682));
    LocalMux I__1467 (
            .O(N__8682),
            .I(\d4.trans_up_1_11 ));
    CascadeMux I__1466 (
            .O(N__8679),
            .I(\d4.trans_up_1_13_cascade_ ));
    InMux I__1465 (
            .O(N__8676),
            .I(N__8673));
    LocalMux I__1464 (
            .O(N__8673),
            .I(\d4.trans_up_1_10 ));
    CascadeMux I__1463 (
            .O(N__8670),
            .I(\d1.g2Z0Z_1_cascade_ ));
    CascadeMux I__1462 (
            .O(N__8667),
            .I(\d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_ ));
    InMux I__1461 (
            .O(N__8664),
            .I(N__8659));
    CascadeMux I__1460 (
            .O(N__8663),
            .I(N__8656));
    InMux I__1459 (
            .O(N__8662),
            .I(N__8652));
    LocalMux I__1458 (
            .O(N__8659),
            .I(N__8649));
    InMux I__1457 (
            .O(N__8656),
            .I(N__8646));
    InMux I__1456 (
            .O(N__8655),
            .I(N__8643));
    LocalMux I__1455 (
            .O(N__8652),
            .I(N__8640));
    Span4Mux_v I__1454 (
            .O(N__8649),
            .I(N__8635));
    LocalMux I__1453 (
            .O(N__8646),
            .I(N__8635));
    LocalMux I__1452 (
            .O(N__8643),
            .I(\a.countZ0Z_0 ));
    Odrv4 I__1451 (
            .O(N__8640),
            .I(\a.countZ0Z_0 ));
    Odrv4 I__1450 (
            .O(N__8635),
            .I(\a.countZ0Z_0 ));
    InMux I__1449 (
            .O(N__8628),
            .I(N__8625));
    LocalMux I__1448 (
            .O(N__8625),
            .I(N__8622));
    Odrv4 I__1447 (
            .O(N__8622),
            .I(\d3.trans_up_1_15_1 ));
    CascadeMux I__1446 (
            .O(N__8619),
            .I(N__8616));
    InMux I__1445 (
            .O(N__8616),
            .I(N__8613));
    LocalMux I__1444 (
            .O(N__8613),
            .I(N__8607));
    InMux I__1443 (
            .O(N__8612),
            .I(N__8604));
    InMux I__1442 (
            .O(N__8611),
            .I(N__8601));
    InMux I__1441 (
            .O(N__8610),
            .I(N__8598));
    Span4Mux_h I__1440 (
            .O(N__8607),
            .I(N__8595));
    LocalMux I__1439 (
            .O(N__8604),
            .I(N__8592));
    LocalMux I__1438 (
            .O(N__8601),
            .I(N__8589));
    LocalMux I__1437 (
            .O(N__8598),
            .I(\d1.countZ0Z_12 ));
    Odrv4 I__1436 (
            .O(N__8595),
            .I(\d1.countZ0Z_12 ));
    Odrv4 I__1435 (
            .O(N__8592),
            .I(\d1.countZ0Z_12 ));
    Odrv4 I__1434 (
            .O(N__8589),
            .I(\d1.countZ0Z_12 ));
    InMux I__1433 (
            .O(N__8580),
            .I(N__8577));
    LocalMux I__1432 (
            .O(N__8577),
            .I(N__8574));
    Span4Mux_v I__1431 (
            .O(N__8574),
            .I(N__8571));
    Sp12to4 I__1430 (
            .O(N__8571),
            .I(N__8568));
    Span12Mux_h I__1429 (
            .O(N__8568),
            .I(N__8565));
    Odrv12 I__1428 (
            .O(N__8565),
            .I(switch_cancel_c));
    InMux I__1427 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__1426 (
            .O(N__8559),
            .I(N__8556));
    Span4Mux_v I__1425 (
            .O(N__8556),
            .I(N__8553));
    Odrv4 I__1424 (
            .O(N__8553),
            .I(\d3.syncZ0Z_0 ));
    InMux I__1423 (
            .O(N__8550),
            .I(N__8547));
    LocalMux I__1422 (
            .O(N__8547),
            .I(N__8544));
    Odrv12 I__1421 (
            .O(N__8544),
            .I(\d1.g2_7_1 ));
    InMux I__1420 (
            .O(N__8541),
            .I(N__8538));
    LocalMux I__1419 (
            .O(N__8538),
            .I(N__8535));
    Span4Mux_h I__1418 (
            .O(N__8535),
            .I(N__8532));
    Odrv4 I__1417 (
            .O(N__8532),
            .I(\d2.syncZ0Z_0 ));
    IoInMux I__1416 (
            .O(N__8529),
            .I(N__8526));
    LocalMux I__1415 (
            .O(N__8526),
            .I(N__8523));
    IoSpan4Mux I__1414 (
            .O(N__8523),
            .I(N__8520));
    Span4Mux_s2_v I__1413 (
            .O(N__8520),
            .I(N__8517));
    Span4Mux_v I__1412 (
            .O(N__8517),
            .I(N__8514));
    Span4Mux_v I__1411 (
            .O(N__8514),
            .I(N__8511));
    Odrv4 I__1410 (
            .O(N__8511),
            .I(\d4.idle_i ));
    InMux I__1409 (
            .O(N__8508),
            .I(N__8505));
    LocalMux I__1408 (
            .O(N__8505),
            .I(\d1.g2_12_0 ));
    CascadeMux I__1407 (
            .O(N__8502),
            .I(\d1.g2Z0Z_12_cascade_ ));
    InMux I__1406 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__1405 (
            .O(N__8496),
            .I(N__8492));
    InMux I__1404 (
            .O(N__8495),
            .I(N__8489));
    Span4Mux_h I__1403 (
            .O(N__8492),
            .I(N__8486));
    LocalMux I__1402 (
            .O(N__8489),
            .I(prescalerZ0Z_10));
    Odrv4 I__1401 (
            .O(N__8486),
            .I(prescalerZ0Z_10));
    InMux I__1400 (
            .O(N__8481),
            .I(N__8477));
    InMux I__1399 (
            .O(N__8480),
            .I(N__8474));
    LocalMux I__1398 (
            .O(N__8477),
            .I(prescalerZ0Z_11));
    LocalMux I__1397 (
            .O(N__8474),
            .I(prescalerZ0Z_11));
    CascadeMux I__1396 (
            .O(N__8469),
            .I(N__8465));
    InMux I__1395 (
            .O(N__8468),
            .I(N__8462));
    InMux I__1394 (
            .O(N__8465),
            .I(N__8459));
    LocalMux I__1393 (
            .O(N__8462),
            .I(prescalerZ0Z_9));
    LocalMux I__1392 (
            .O(N__8459),
            .I(prescalerZ0Z_9));
    InMux I__1391 (
            .O(N__8454),
            .I(N__8450));
    InMux I__1390 (
            .O(N__8453),
            .I(N__8447));
    LocalMux I__1389 (
            .O(N__8450),
            .I(prescalerZ0Z_12));
    LocalMux I__1388 (
            .O(N__8447),
            .I(prescalerZ0Z_12));
    CascadeMux I__1387 (
            .O(N__8442),
            .I(N__8439));
    InMux I__1386 (
            .O(N__8439),
            .I(N__8436));
    LocalMux I__1385 (
            .O(N__8436),
            .I(N__8433));
    Span4Mux_h I__1384 (
            .O(N__8433),
            .I(N__8430));
    Odrv4 I__1383 (
            .O(N__8430),
            .I(decrement_time_0_prescaler10_5_and));
    InMux I__1382 (
            .O(N__8427),
            .I(N__8423));
    InMux I__1381 (
            .O(N__8426),
            .I(N__8420));
    LocalMux I__1380 (
            .O(N__8423),
            .I(N__8417));
    LocalMux I__1379 (
            .O(N__8420),
            .I(prescalerZ0Z_25));
    Odrv4 I__1378 (
            .O(N__8417),
            .I(prescalerZ0Z_25));
    InMux I__1377 (
            .O(N__8412),
            .I(N__8408));
    InMux I__1376 (
            .O(N__8411),
            .I(N__8405));
    LocalMux I__1375 (
            .O(N__8408),
            .I(prescalerZ0Z_27));
    LocalMux I__1374 (
            .O(N__8405),
            .I(prescalerZ0Z_27));
    CascadeMux I__1373 (
            .O(N__8400),
            .I(N__8396));
    InMux I__1372 (
            .O(N__8399),
            .I(N__8393));
    InMux I__1371 (
            .O(N__8396),
            .I(N__8390));
    LocalMux I__1370 (
            .O(N__8393),
            .I(prescalerZ0Z_17));
    LocalMux I__1369 (
            .O(N__8390),
            .I(prescalerZ0Z_17));
    InMux I__1368 (
            .O(N__8385),
            .I(N__8381));
    InMux I__1367 (
            .O(N__8384),
            .I(N__8378));
    LocalMux I__1366 (
            .O(N__8381),
            .I(prescalerZ0Z_19));
    LocalMux I__1365 (
            .O(N__8378),
            .I(prescalerZ0Z_19));
    CascadeMux I__1364 (
            .O(N__8373),
            .I(N__8370));
    InMux I__1363 (
            .O(N__8370),
            .I(N__8367));
    LocalMux I__1362 (
            .O(N__8367),
            .I(N__8364));
    Span4Mux_h I__1361 (
            .O(N__8364),
            .I(N__8361));
    Odrv4 I__1360 (
            .O(N__8361),
            .I(decrement_time_0_prescaler10_6_and));
    CascadeMux I__1359 (
            .O(N__8358),
            .I(\d1.g2_7_2_cascade_ ));
    CascadeMux I__1358 (
            .O(N__8355),
            .I(\d1.mins27_1_cascade_ ));
    CascadeMux I__1357 (
            .O(N__8352),
            .I(\d1.g2Z0Z_0_cascade_ ));
    InMux I__1356 (
            .O(N__8349),
            .I(N__8346));
    LocalMux I__1355 (
            .O(N__8346),
            .I(N__8343));
    Odrv4 I__1354 (
            .O(N__8343),
            .I(\d1.g0_1_a5_0_9 ));
    InMux I__1353 (
            .O(N__8340),
            .I(N__8337));
    LocalMux I__1352 (
            .O(N__8337),
            .I(N__8334));
    Odrv4 I__1351 (
            .O(N__8334),
            .I(\d1.g0_1_a5_0_8 ));
    InMux I__1350 (
            .O(N__8331),
            .I(N__8328));
    LocalMux I__1349 (
            .O(N__8328),
            .I(N__8325));
    Odrv12 I__1348 (
            .O(N__8325),
            .I(\d1.g0_0_0_a4_2_0 ));
    InMux I__1347 (
            .O(N__8322),
            .I(N__8319));
    LocalMux I__1346 (
            .O(N__8319),
            .I(\d1.gZ0Z2 ));
    InMux I__1345 (
            .O(N__8316),
            .I(N__8310));
    InMux I__1344 (
            .O(N__8315),
            .I(N__8310));
    LocalMux I__1343 (
            .O(N__8310),
            .I(N__8305));
    InMux I__1342 (
            .O(N__8309),
            .I(N__8300));
    InMux I__1341 (
            .O(N__8308),
            .I(N__8297));
    Span4Mux_h I__1340 (
            .O(N__8305),
            .I(N__8294));
    InMux I__1339 (
            .O(N__8304),
            .I(N__8289));
    InMux I__1338 (
            .O(N__8303),
            .I(N__8289));
    LocalMux I__1337 (
            .O(N__8300),
            .I(\d1.countZ0Z_0 ));
    LocalMux I__1336 (
            .O(N__8297),
            .I(\d1.countZ0Z_0 ));
    Odrv4 I__1335 (
            .O(N__8294),
            .I(\d1.countZ0Z_0 ));
    LocalMux I__1334 (
            .O(N__8289),
            .I(\d1.countZ0Z_0 ));
    CascadeMux I__1333 (
            .O(N__8280),
            .I(N__8277));
    InMux I__1332 (
            .O(N__8277),
            .I(N__8271));
    InMux I__1331 (
            .O(N__8276),
            .I(N__8271));
    LocalMux I__1330 (
            .O(N__8271),
            .I(N__8266));
    InMux I__1329 (
            .O(N__8270),
            .I(N__8263));
    InMux I__1328 (
            .O(N__8269),
            .I(N__8260));
    Span4Mux_h I__1327 (
            .O(N__8266),
            .I(N__8257));
    LocalMux I__1326 (
            .O(N__8263),
            .I(N__8254));
    LocalMux I__1325 (
            .O(N__8260),
            .I(\d1.countZ0Z_11 ));
    Odrv4 I__1324 (
            .O(N__8257),
            .I(\d1.countZ0Z_11 ));
    Odrv4 I__1323 (
            .O(N__8254),
            .I(\d1.countZ0Z_11 ));
    CascadeMux I__1322 (
            .O(N__8247),
            .I(N__8244));
    InMux I__1321 (
            .O(N__8244),
            .I(N__8241));
    LocalMux I__1320 (
            .O(N__8241),
            .I(decrement_time_0_prescaler10_2_and));
    CascadeMux I__1319 (
            .O(N__8238),
            .I(N__8235));
    InMux I__1318 (
            .O(N__8235),
            .I(N__8232));
    LocalMux I__1317 (
            .O(N__8232),
            .I(decrement_time_0_prescaler10_3_and));
    CascadeMux I__1316 (
            .O(N__8229),
            .I(N__8226));
    InMux I__1315 (
            .O(N__8226),
            .I(N__8223));
    LocalMux I__1314 (
            .O(N__8223),
            .I(N__8220));
    Odrv4 I__1313 (
            .O(N__8220),
            .I(decrement_time_0_prescaler10_4_and));
    InMux I__1312 (
            .O(N__8217),
            .I(decrement_time_0_prescaler10));
    InMux I__1311 (
            .O(N__8214),
            .I(N__8211));
    LocalMux I__1310 (
            .O(N__8211),
            .I(N__8208));
    Span4Mux_h I__1309 (
            .O(N__8208),
            .I(N__8205));
    Odrv4 I__1308 (
            .O(N__8205),
            .I(prescaler_1_cry_12_THRU_CO));
    InMux I__1307 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1306 (
            .O(N__8199),
            .I(N__8194));
    CascadeMux I__1305 (
            .O(N__8198),
            .I(N__8191));
    InMux I__1304 (
            .O(N__8197),
            .I(N__8188));
    Span4Mux_v I__1303 (
            .O(N__8194),
            .I(N__8185));
    InMux I__1302 (
            .O(N__8191),
            .I(N__8182));
    LocalMux I__1301 (
            .O(N__8188),
            .I(prescalerZ0Z_13));
    Odrv4 I__1300 (
            .O(N__8185),
            .I(prescalerZ0Z_13));
    LocalMux I__1299 (
            .O(N__8182),
            .I(prescalerZ0Z_13));
    InMux I__1298 (
            .O(N__8175),
            .I(N__8172));
    LocalMux I__1297 (
            .O(N__8172),
            .I(N__8169));
    Span4Mux_v I__1296 (
            .O(N__8169),
            .I(N__8166));
    Odrv4 I__1295 (
            .O(N__8166),
            .I(prescaler_1_cry_13_THRU_CO));
    InMux I__1294 (
            .O(N__8163),
            .I(N__8160));
    LocalMux I__1293 (
            .O(N__8160),
            .I(N__8157));
    Span4Mux_v I__1292 (
            .O(N__8157),
            .I(N__8152));
    InMux I__1291 (
            .O(N__8156),
            .I(N__8147));
    InMux I__1290 (
            .O(N__8155),
            .I(N__8147));
    Odrv4 I__1289 (
            .O(N__8152),
            .I(prescalerZ0Z_14));
    LocalMux I__1288 (
            .O(N__8147),
            .I(prescalerZ0Z_14));
    InMux I__1287 (
            .O(N__8142),
            .I(N__8139));
    LocalMux I__1286 (
            .O(N__8139),
            .I(N__8136));
    Span4Mux_h I__1285 (
            .O(N__8136),
            .I(N__8133));
    Span4Mux_v I__1284 (
            .O(N__8133),
            .I(N__8130));
    Odrv4 I__1283 (
            .O(N__8130),
            .I(prescaler_1_cry_14_THRU_CO));
    InMux I__1282 (
            .O(N__8127),
            .I(N__8124));
    LocalMux I__1281 (
            .O(N__8124),
            .I(N__8121));
    Span4Mux_v I__1280 (
            .O(N__8121),
            .I(N__8116));
    InMux I__1279 (
            .O(N__8120),
            .I(N__8111));
    InMux I__1278 (
            .O(N__8119),
            .I(N__8111));
    Odrv4 I__1277 (
            .O(N__8116),
            .I(prescalerZ0Z_15));
    LocalMux I__1276 (
            .O(N__8111),
            .I(prescalerZ0Z_15));
    InMux I__1275 (
            .O(N__8106),
            .I(N__8103));
    LocalMux I__1274 (
            .O(N__8103),
            .I(N__8100));
    Span4Mux_v I__1273 (
            .O(N__8100),
            .I(N__8097));
    Odrv4 I__1272 (
            .O(N__8097),
            .I(prescaler_1_cry_15_THRU_CO));
    InMux I__1271 (
            .O(N__8094),
            .I(N__8091));
    LocalMux I__1270 (
            .O(N__8091),
            .I(N__8087));
    CascadeMux I__1269 (
            .O(N__8090),
            .I(N__8084));
    Span4Mux_v I__1268 (
            .O(N__8087),
            .I(N__8080));
    InMux I__1267 (
            .O(N__8084),
            .I(N__8075));
    InMux I__1266 (
            .O(N__8083),
            .I(N__8075));
    Odrv4 I__1265 (
            .O(N__8080),
            .I(prescalerZ0Z_16));
    LocalMux I__1264 (
            .O(N__8075),
            .I(prescalerZ0Z_16));
    InMux I__1263 (
            .O(N__8070),
            .I(N__8067));
    LocalMux I__1262 (
            .O(N__8067),
            .I(N__8064));
    Span4Mux_v I__1261 (
            .O(N__8064),
            .I(N__8061));
    Odrv4 I__1260 (
            .O(N__8061),
            .I(prescaler_1_cry_17_THRU_CO));
    CEMux I__1259 (
            .O(N__8058),
            .I(N__8037));
    CEMux I__1258 (
            .O(N__8057),
            .I(N__8037));
    CEMux I__1257 (
            .O(N__8056),
            .I(N__8037));
    CEMux I__1256 (
            .O(N__8055),
            .I(N__8037));
    CEMux I__1255 (
            .O(N__8054),
            .I(N__8037));
    CEMux I__1254 (
            .O(N__8053),
            .I(N__8037));
    CEMux I__1253 (
            .O(N__8052),
            .I(N__8037));
    GlobalMux I__1252 (
            .O(N__8037),
            .I(N__8034));
    gio2CtrlBuf I__1251 (
            .O(N__8034),
            .I(un1_state_3_g));
    InMux I__1250 (
            .O(N__8031),
            .I(N__8028));
    LocalMux I__1249 (
            .O(N__8028),
            .I(N__8024));
    InMux I__1248 (
            .O(N__8027),
            .I(N__8020));
    Span4Mux_v I__1247 (
            .O(N__8024),
            .I(N__8017));
    InMux I__1246 (
            .O(N__8023),
            .I(N__8014));
    LocalMux I__1245 (
            .O(N__8020),
            .I(prescalerZ0Z_20));
    Odrv4 I__1244 (
            .O(N__8017),
            .I(prescalerZ0Z_20));
    LocalMux I__1243 (
            .O(N__8014),
            .I(prescalerZ0Z_20));
    InMux I__1242 (
            .O(N__8007),
            .I(N__8004));
    LocalMux I__1241 (
            .O(N__8004),
            .I(N__8000));
    InMux I__1240 (
            .O(N__8003),
            .I(N__7996));
    Span4Mux_v I__1239 (
            .O(N__8000),
            .I(N__7993));
    InMux I__1238 (
            .O(N__7999),
            .I(N__7990));
    LocalMux I__1237 (
            .O(N__7996),
            .I(prescalerZ0Z_21));
    Odrv4 I__1236 (
            .O(N__7993),
            .I(prescalerZ0Z_21));
    LocalMux I__1235 (
            .O(N__7990),
            .I(prescalerZ0Z_21));
    CascadeMux I__1234 (
            .O(N__7983),
            .I(N__7980));
    InMux I__1233 (
            .O(N__7980),
            .I(N__7976));
    CascadeMux I__1232 (
            .O(N__7979),
            .I(N__7973));
    LocalMux I__1231 (
            .O(N__7976),
            .I(N__7969));
    InMux I__1230 (
            .O(N__7973),
            .I(N__7966));
    InMux I__1229 (
            .O(N__7972),
            .I(N__7963));
    Span4Mux_v I__1228 (
            .O(N__7969),
            .I(N__7958));
    LocalMux I__1227 (
            .O(N__7966),
            .I(N__7958));
    LocalMux I__1226 (
            .O(N__7963),
            .I(prescalerZ0Z_22));
    Odrv4 I__1225 (
            .O(N__7958),
            .I(prescalerZ0Z_22));
    InMux I__1224 (
            .O(N__7953),
            .I(N__7950));
    LocalMux I__1223 (
            .O(N__7950),
            .I(N__7947));
    Span4Mux_v I__1222 (
            .O(N__7947),
            .I(N__7942));
    InMux I__1221 (
            .O(N__7946),
            .I(N__7937));
    InMux I__1220 (
            .O(N__7945),
            .I(N__7937));
    Odrv4 I__1219 (
            .O(N__7942),
            .I(prescalerZ0Z_18));
    LocalMux I__1218 (
            .O(N__7937),
            .I(prescalerZ0Z_18));
    CascadeMux I__1217 (
            .O(N__7932),
            .I(N__7929));
    InMux I__1216 (
            .O(N__7929),
            .I(N__7926));
    LocalMux I__1215 (
            .O(N__7926),
            .I(decrement_time_0_prescaler10_0_and));
    CascadeMux I__1214 (
            .O(N__7923),
            .I(N__7920));
    InMux I__1213 (
            .O(N__7920),
            .I(N__7917));
    LocalMux I__1212 (
            .O(N__7917),
            .I(decrement_time_0_prescaler10_1_and));
    InMux I__1211 (
            .O(N__7914),
            .I(N__7911));
    LocalMux I__1210 (
            .O(N__7911),
            .I(N__7908));
    Span12Mux_v I__1209 (
            .O(N__7908),
            .I(N__7905));
    Odrv12 I__1208 (
            .O(N__7905),
            .I(prescaler_1_cry_7_THRU_CO));
    InMux I__1207 (
            .O(N__7902),
            .I(N__7898));
    InMux I__1206 (
            .O(N__7901),
            .I(N__7895));
    LocalMux I__1205 (
            .O(N__7898),
            .I(N__7892));
    LocalMux I__1204 (
            .O(N__7895),
            .I(N__7886));
    Span4Mux_v I__1203 (
            .O(N__7892),
            .I(N__7886));
    InMux I__1202 (
            .O(N__7891),
            .I(N__7883));
    Odrv4 I__1201 (
            .O(N__7886),
            .I(prescalerZ0Z_8));
    LocalMux I__1200 (
            .O(N__7883),
            .I(prescalerZ0Z_8));
    InMux I__1199 (
            .O(N__7878),
            .I(N__7875));
    LocalMux I__1198 (
            .O(N__7875),
            .I(N__7872));
    Span4Mux_v I__1197 (
            .O(N__7872),
            .I(N__7869));
    Odrv4 I__1196 (
            .O(N__7869),
            .I(prescaler_1_cry_22_THRU_CO));
    InMux I__1195 (
            .O(N__7866),
            .I(N__7863));
    LocalMux I__1194 (
            .O(N__7863),
            .I(N__7860));
    Span4Mux_v I__1193 (
            .O(N__7860),
            .I(N__7855));
    InMux I__1192 (
            .O(N__7859),
            .I(N__7850));
    InMux I__1191 (
            .O(N__7858),
            .I(N__7850));
    Odrv4 I__1190 (
            .O(N__7855),
            .I(prescalerZ0Z_23));
    LocalMux I__1189 (
            .O(N__7850),
            .I(prescalerZ0Z_23));
    InMux I__1188 (
            .O(N__7845),
            .I(N__7842));
    LocalMux I__1187 (
            .O(N__7842),
            .I(N__7839));
    Span4Mux_v I__1186 (
            .O(N__7839),
            .I(N__7836));
    Odrv4 I__1185 (
            .O(N__7836),
            .I(prescaler_1_cry_23_THRU_CO));
    InMux I__1184 (
            .O(N__7833),
            .I(N__7830));
    LocalMux I__1183 (
            .O(N__7830),
            .I(N__7825));
    CascadeMux I__1182 (
            .O(N__7829),
            .I(N__7822));
    InMux I__1181 (
            .O(N__7828),
            .I(N__7819));
    Sp12to4 I__1180 (
            .O(N__7825),
            .I(N__7816));
    InMux I__1179 (
            .O(N__7822),
            .I(N__7813));
    LocalMux I__1178 (
            .O(N__7819),
            .I(prescalerZ0Z_24));
    Odrv12 I__1177 (
            .O(N__7816),
            .I(prescalerZ0Z_24));
    LocalMux I__1176 (
            .O(N__7813),
            .I(prescalerZ0Z_24));
    InMux I__1175 (
            .O(N__7806),
            .I(N__7803));
    LocalMux I__1174 (
            .O(N__7803),
            .I(N__7800));
    Span4Mux_h I__1173 (
            .O(N__7800),
            .I(N__7797));
    Span4Mux_v I__1172 (
            .O(N__7797),
            .I(N__7794));
    Odrv4 I__1171 (
            .O(N__7794),
            .I(prescaler_1_cry_25_THRU_CO));
    InMux I__1170 (
            .O(N__7791),
            .I(N__7788));
    LocalMux I__1169 (
            .O(N__7788),
            .I(N__7785));
    Span4Mux_v I__1168 (
            .O(N__7785),
            .I(N__7780));
    InMux I__1167 (
            .O(N__7784),
            .I(N__7775));
    InMux I__1166 (
            .O(N__7783),
            .I(N__7775));
    Odrv4 I__1165 (
            .O(N__7780),
            .I(prescalerZ0Z_26));
    LocalMux I__1164 (
            .O(N__7775),
            .I(prescalerZ0Z_26));
    InMux I__1163 (
            .O(N__7770),
            .I(N__7767));
    LocalMux I__1162 (
            .O(N__7767),
            .I(N__7764));
    Span4Mux_v I__1161 (
            .O(N__7764),
            .I(N__7761));
    Span4Mux_v I__1160 (
            .O(N__7761),
            .I(N__7758));
    Odrv4 I__1159 (
            .O(N__7758),
            .I(prescaler_1_cry_19_THRU_CO));
    InMux I__1158 (
            .O(N__7755),
            .I(N__7752));
    LocalMux I__1157 (
            .O(N__7752),
            .I(N__7749));
    Span4Mux_v I__1156 (
            .O(N__7749),
            .I(N__7746));
    Odrv4 I__1155 (
            .O(N__7746),
            .I(prescaler_1_cry_20_THRU_CO));
    InMux I__1154 (
            .O(N__7743),
            .I(N__7740));
    LocalMux I__1153 (
            .O(N__7740),
            .I(N__7737));
    Span4Mux_v I__1152 (
            .O(N__7737),
            .I(N__7734));
    Odrv4 I__1151 (
            .O(N__7734),
            .I(prescaler_1_cry_21_THRU_CO));
    InMux I__1150 (
            .O(N__7731),
            .I(prescaler_1_cry_18));
    InMux I__1149 (
            .O(N__7728),
            .I(prescaler_1_cry_19));
    InMux I__1148 (
            .O(N__7725),
            .I(prescaler_1_cry_20));
    InMux I__1147 (
            .O(N__7722),
            .I(prescaler_1_cry_21));
    InMux I__1146 (
            .O(N__7719),
            .I(prescaler_1_cry_22));
    InMux I__1145 (
            .O(N__7716),
            .I(prescaler_1_cry_23));
    InMux I__1144 (
            .O(N__7713),
            .I(bfn_8_18_0_));
    InMux I__1143 (
            .O(N__7710),
            .I(prescaler_1_cry_25));
    InMux I__1142 (
            .O(N__7707),
            .I(prescaler_1_cry_26));
    InMux I__1141 (
            .O(N__7704),
            .I(prescaler_1_cry_9));
    InMux I__1140 (
            .O(N__7701),
            .I(prescaler_1_cry_10));
    InMux I__1139 (
            .O(N__7698),
            .I(prescaler_1_cry_11));
    InMux I__1138 (
            .O(N__7695),
            .I(prescaler_1_cry_12));
    InMux I__1137 (
            .O(N__7692),
            .I(prescaler_1_cry_13));
    InMux I__1136 (
            .O(N__7689),
            .I(prescaler_1_cry_14));
    InMux I__1135 (
            .O(N__7686),
            .I(prescaler_1_cry_15));
    InMux I__1134 (
            .O(N__7683),
            .I(bfn_8_17_0_));
    InMux I__1133 (
            .O(N__7680),
            .I(prescaler_1_cry_17));
    CascadeMux I__1132 (
            .O(N__7677),
            .I(N__7671));
    InMux I__1131 (
            .O(N__7676),
            .I(N__7666));
    InMux I__1130 (
            .O(N__7675),
            .I(N__7666));
    InMux I__1129 (
            .O(N__7674),
            .I(N__7663));
    InMux I__1128 (
            .O(N__7671),
            .I(N__7660));
    LocalMux I__1127 (
            .O(N__7666),
            .I(prescalerZ0Z_0));
    LocalMux I__1126 (
            .O(N__7663),
            .I(prescalerZ0Z_0));
    LocalMux I__1125 (
            .O(N__7660),
            .I(prescalerZ0Z_0));
    CascadeMux I__1124 (
            .O(N__7653),
            .I(N__7649));
    InMux I__1123 (
            .O(N__7652),
            .I(N__7645));
    InMux I__1122 (
            .O(N__7649),
            .I(N__7642));
    InMux I__1121 (
            .O(N__7648),
            .I(N__7639));
    LocalMux I__1120 (
            .O(N__7645),
            .I(prescalerZ0Z_1));
    LocalMux I__1119 (
            .O(N__7642),
            .I(prescalerZ0Z_1));
    LocalMux I__1118 (
            .O(N__7639),
            .I(prescalerZ0Z_1));
    InMux I__1117 (
            .O(N__7632),
            .I(N__7628));
    InMux I__1116 (
            .O(N__7631),
            .I(N__7625));
    LocalMux I__1115 (
            .O(N__7628),
            .I(N__7622));
    LocalMux I__1114 (
            .O(N__7625),
            .I(prescalerZ0Z_2));
    Odrv4 I__1113 (
            .O(N__7622),
            .I(prescalerZ0Z_2));
    InMux I__1112 (
            .O(N__7617),
            .I(prescaler_1_cry_1));
    InMux I__1111 (
            .O(N__7614),
            .I(N__7610));
    InMux I__1110 (
            .O(N__7613),
            .I(N__7607));
    LocalMux I__1109 (
            .O(N__7610),
            .I(N__7604));
    LocalMux I__1108 (
            .O(N__7607),
            .I(prescalerZ0Z_3));
    Odrv4 I__1107 (
            .O(N__7604),
            .I(prescalerZ0Z_3));
    InMux I__1106 (
            .O(N__7599),
            .I(prescaler_1_cry_2));
    InMux I__1105 (
            .O(N__7596),
            .I(N__7592));
    InMux I__1104 (
            .O(N__7595),
            .I(N__7589));
    LocalMux I__1103 (
            .O(N__7592),
            .I(prescalerZ0Z_4));
    LocalMux I__1102 (
            .O(N__7589),
            .I(prescalerZ0Z_4));
    InMux I__1101 (
            .O(N__7584),
            .I(prescaler_1_cry_3));
    CascadeMux I__1100 (
            .O(N__7581),
            .I(N__7577));
    InMux I__1099 (
            .O(N__7580),
            .I(N__7574));
    InMux I__1098 (
            .O(N__7577),
            .I(N__7571));
    LocalMux I__1097 (
            .O(N__7574),
            .I(prescalerZ0Z_5));
    LocalMux I__1096 (
            .O(N__7571),
            .I(prescalerZ0Z_5));
    InMux I__1095 (
            .O(N__7566),
            .I(prescaler_1_cry_4));
    InMux I__1094 (
            .O(N__7563),
            .I(N__7559));
    InMux I__1093 (
            .O(N__7562),
            .I(N__7556));
    LocalMux I__1092 (
            .O(N__7559),
            .I(prescalerZ0Z_6));
    LocalMux I__1091 (
            .O(N__7556),
            .I(prescalerZ0Z_6));
    InMux I__1090 (
            .O(N__7551),
            .I(prescaler_1_cry_5));
    InMux I__1089 (
            .O(N__7548),
            .I(N__7544));
    InMux I__1088 (
            .O(N__7547),
            .I(N__7541));
    LocalMux I__1087 (
            .O(N__7544),
            .I(prescalerZ0Z_7));
    LocalMux I__1086 (
            .O(N__7541),
            .I(prescalerZ0Z_7));
    InMux I__1085 (
            .O(N__7536),
            .I(prescaler_1_cry_6));
    InMux I__1084 (
            .O(N__7533),
            .I(prescaler_1_cry_7));
    InMux I__1083 (
            .O(N__7530),
            .I(bfn_8_16_0_));
    InMux I__1082 (
            .O(N__7527),
            .I(\a.count_1_cry_20 ));
    InMux I__1081 (
            .O(N__7524),
            .I(N__7520));
    InMux I__1080 (
            .O(N__7523),
            .I(N__7517));
    LocalMux I__1079 (
            .O(N__7520),
            .I(N__7514));
    LocalMux I__1078 (
            .O(N__7517),
            .I(\a.countZ0Z_22 ));
    Odrv4 I__1077 (
            .O(N__7514),
            .I(\a.countZ0Z_22 ));
    InMux I__1076 (
            .O(N__7509),
            .I(\a.count_1_cry_21 ));
    InMux I__1075 (
            .O(N__7506),
            .I(N__7502));
    InMux I__1074 (
            .O(N__7505),
            .I(N__7499));
    LocalMux I__1073 (
            .O(N__7502),
            .I(\a.countZ0Z_23 ));
    LocalMux I__1072 (
            .O(N__7499),
            .I(\a.countZ0Z_23 ));
    InMux I__1071 (
            .O(N__7494),
            .I(\a.count_1_cry_22 ));
    InMux I__1070 (
            .O(N__7491),
            .I(N__7487));
    InMux I__1069 (
            .O(N__7490),
            .I(N__7484));
    LocalMux I__1068 (
            .O(N__7487),
            .I(\a.countZ0Z_24 ));
    LocalMux I__1067 (
            .O(N__7484),
            .I(\a.countZ0Z_24 ));
    InMux I__1066 (
            .O(N__7479),
            .I(\a.count_1_cry_23 ));
    InMux I__1065 (
            .O(N__7476),
            .I(bfn_8_14_0_));
    CascadeMux I__1064 (
            .O(N__7473),
            .I(N__7469));
    InMux I__1063 (
            .O(N__7472),
            .I(N__7466));
    InMux I__1062 (
            .O(N__7469),
            .I(N__7463));
    LocalMux I__1061 (
            .O(N__7466),
            .I(\a.countZ0Z_25 ));
    LocalMux I__1060 (
            .O(N__7463),
            .I(\a.countZ0Z_25 ));
    InMux I__1059 (
            .O(N__7458),
            .I(N__7454));
    InMux I__1058 (
            .O(N__7457),
            .I(N__7451));
    LocalMux I__1057 (
            .O(N__7454),
            .I(\a.countZ0Z_18 ));
    LocalMux I__1056 (
            .O(N__7451),
            .I(\a.countZ0Z_18 ));
    InMux I__1055 (
            .O(N__7446),
            .I(N__7442));
    InMux I__1054 (
            .O(N__7445),
            .I(N__7439));
    LocalMux I__1053 (
            .O(N__7442),
            .I(N__7436));
    LocalMux I__1052 (
            .O(N__7439),
            .I(\a.countZ0Z_21 ));
    Odrv4 I__1051 (
            .O(N__7436),
            .I(\a.countZ0Z_21 ));
    CascadeMux I__1050 (
            .O(N__7431),
            .I(N__7427));
    InMux I__1049 (
            .O(N__7430),
            .I(N__7424));
    InMux I__1048 (
            .O(N__7427),
            .I(N__7421));
    LocalMux I__1047 (
            .O(N__7424),
            .I(\a.countZ0Z_20 ));
    LocalMux I__1046 (
            .O(N__7421),
            .I(\a.countZ0Z_20 ));
    InMux I__1045 (
            .O(N__7416),
            .I(N__7412));
    InMux I__1044 (
            .O(N__7415),
            .I(N__7409));
    LocalMux I__1043 (
            .O(N__7412),
            .I(\a.countZ0Z_19 ));
    LocalMux I__1042 (
            .O(N__7409),
            .I(\a.countZ0Z_19 ));
    InMux I__1041 (
            .O(N__7404),
            .I(N__7401));
    LocalMux I__1040 (
            .O(N__7401),
            .I(\a.BUZZER3_15 ));
    InMux I__1039 (
            .O(N__7398),
            .I(N__7394));
    InMux I__1038 (
            .O(N__7397),
            .I(N__7391));
    LocalMux I__1037 (
            .O(N__7394),
            .I(\a.countZ0Z_12 ));
    LocalMux I__1036 (
            .O(N__7391),
            .I(\a.countZ0Z_12 ));
    InMux I__1035 (
            .O(N__7386),
            .I(N__7383));
    LocalMux I__1034 (
            .O(N__7383),
            .I(\a.count_1_12 ));
    InMux I__1033 (
            .O(N__7380),
            .I(\a.count_1_cry_11 ));
    InMux I__1032 (
            .O(N__7377),
            .I(N__7373));
    InMux I__1031 (
            .O(N__7376),
            .I(N__7370));
    LocalMux I__1030 (
            .O(N__7373),
            .I(\a.countZ0Z_13 ));
    LocalMux I__1029 (
            .O(N__7370),
            .I(\a.countZ0Z_13 ));
    InMux I__1028 (
            .O(N__7365),
            .I(N__7362));
    LocalMux I__1027 (
            .O(N__7362),
            .I(\a.count_1_13 ));
    InMux I__1026 (
            .O(N__7359),
            .I(\a.count_1_cry_12 ));
    InMux I__1025 (
            .O(N__7356),
            .I(N__7352));
    InMux I__1024 (
            .O(N__7355),
            .I(N__7349));
    LocalMux I__1023 (
            .O(N__7352),
            .I(\a.countZ0Z_14 ));
    LocalMux I__1022 (
            .O(N__7349),
            .I(\a.countZ0Z_14 ));
    InMux I__1021 (
            .O(N__7344),
            .I(N__7341));
    LocalMux I__1020 (
            .O(N__7341),
            .I(\a.count_1_14 ));
    InMux I__1019 (
            .O(N__7338),
            .I(\a.count_1_cry_13 ));
    InMux I__1018 (
            .O(N__7335),
            .I(N__7331));
    InMux I__1017 (
            .O(N__7334),
            .I(N__7328));
    LocalMux I__1016 (
            .O(N__7331),
            .I(\a.countZ0Z_15 ));
    LocalMux I__1015 (
            .O(N__7328),
            .I(\a.countZ0Z_15 ));
    InMux I__1014 (
            .O(N__7323),
            .I(\a.count_1_cry_14 ));
    InMux I__1013 (
            .O(N__7320),
            .I(N__7316));
    InMux I__1012 (
            .O(N__7319),
            .I(N__7313));
    LocalMux I__1011 (
            .O(N__7316),
            .I(\a.countZ0Z_16 ));
    LocalMux I__1010 (
            .O(N__7313),
            .I(\a.countZ0Z_16 ));
    InMux I__1009 (
            .O(N__7308),
            .I(\a.count_1_cry_15 ));
    InMux I__1008 (
            .O(N__7305),
            .I(N__7301));
    InMux I__1007 (
            .O(N__7304),
            .I(N__7298));
    LocalMux I__1006 (
            .O(N__7301),
            .I(\a.countZ0Z_17 ));
    LocalMux I__1005 (
            .O(N__7298),
            .I(\a.countZ0Z_17 ));
    InMux I__1004 (
            .O(N__7293),
            .I(bfn_8_13_0_));
    InMux I__1003 (
            .O(N__7290),
            .I(\a.count_1_cry_17 ));
    InMux I__1002 (
            .O(N__7287),
            .I(\a.count_1_cry_18 ));
    InMux I__1001 (
            .O(N__7284),
            .I(\a.count_1_cry_19 ));
    InMux I__1000 (
            .O(N__7281),
            .I(N__7277));
    InMux I__999 (
            .O(N__7280),
            .I(N__7274));
    LocalMux I__998 (
            .O(N__7277),
            .I(\a.countZ0Z_4 ));
    LocalMux I__997 (
            .O(N__7274),
            .I(\a.countZ0Z_4 ));
    InMux I__996 (
            .O(N__7269),
            .I(\a.count_1_cry_3 ));
    InMux I__995 (
            .O(N__7266),
            .I(N__7262));
    InMux I__994 (
            .O(N__7265),
            .I(N__7259));
    LocalMux I__993 (
            .O(N__7262),
            .I(\a.countZ0Z_5 ));
    LocalMux I__992 (
            .O(N__7259),
            .I(\a.countZ0Z_5 ));
    InMux I__991 (
            .O(N__7254),
            .I(\a.count_1_cry_4 ));
    InMux I__990 (
            .O(N__7251),
            .I(N__7247));
    InMux I__989 (
            .O(N__7250),
            .I(N__7244));
    LocalMux I__988 (
            .O(N__7247),
            .I(\a.countZ0Z_6 ));
    LocalMux I__987 (
            .O(N__7244),
            .I(\a.countZ0Z_6 ));
    InMux I__986 (
            .O(N__7239),
            .I(\a.count_1_cry_5 ));
    InMux I__985 (
            .O(N__7236),
            .I(N__7232));
    InMux I__984 (
            .O(N__7235),
            .I(N__7229));
    LocalMux I__983 (
            .O(N__7232),
            .I(\a.countZ0Z_7 ));
    LocalMux I__982 (
            .O(N__7229),
            .I(\a.countZ0Z_7 ));
    InMux I__981 (
            .O(N__7224),
            .I(\a.count_1_cry_6 ));
    CascadeMux I__980 (
            .O(N__7221),
            .I(N__7218));
    InMux I__979 (
            .O(N__7218),
            .I(N__7215));
    LocalMux I__978 (
            .O(N__7215),
            .I(N__7211));
    InMux I__977 (
            .O(N__7214),
            .I(N__7208));
    Odrv4 I__976 (
            .O(N__7211),
            .I(\a.countZ0Z_8 ));
    LocalMux I__975 (
            .O(N__7208),
            .I(\a.countZ0Z_8 ));
    InMux I__974 (
            .O(N__7203),
            .I(N__7200));
    LocalMux I__973 (
            .O(N__7200),
            .I(\a.count_1_8 ));
    InMux I__972 (
            .O(N__7197),
            .I(\a.count_1_cry_7 ));
    InMux I__971 (
            .O(N__7194),
            .I(N__7190));
    InMux I__970 (
            .O(N__7193),
            .I(N__7187));
    LocalMux I__969 (
            .O(N__7190),
            .I(\a.countZ0Z_9 ));
    LocalMux I__968 (
            .O(N__7187),
            .I(\a.countZ0Z_9 ));
    InMux I__967 (
            .O(N__7182),
            .I(bfn_8_12_0_));
    CascadeMux I__966 (
            .O(N__7179),
            .I(N__7176));
    InMux I__965 (
            .O(N__7176),
            .I(N__7172));
    InMux I__964 (
            .O(N__7175),
            .I(N__7169));
    LocalMux I__963 (
            .O(N__7172),
            .I(\a.countZ0Z_10 ));
    LocalMux I__962 (
            .O(N__7169),
            .I(\a.countZ0Z_10 ));
    InMux I__961 (
            .O(N__7164),
            .I(N__7161));
    LocalMux I__960 (
            .O(N__7161),
            .I(\a.count_1_10 ));
    InMux I__959 (
            .O(N__7158),
            .I(\a.count_1_cry_9 ));
    CascadeMux I__958 (
            .O(N__7155),
            .I(N__7152));
    InMux I__957 (
            .O(N__7152),
            .I(N__7148));
    InMux I__956 (
            .O(N__7151),
            .I(N__7145));
    LocalMux I__955 (
            .O(N__7148),
            .I(\a.countZ0Z_11 ));
    LocalMux I__954 (
            .O(N__7145),
            .I(\a.countZ0Z_11 ));
    InMux I__953 (
            .O(N__7140),
            .I(N__7137));
    LocalMux I__952 (
            .O(N__7137),
            .I(\a.count_1_11 ));
    InMux I__951 (
            .O(N__7134),
            .I(\a.count_1_cry_10 ));
    InMux I__950 (
            .O(N__7131),
            .I(N__7127));
    InMux I__949 (
            .O(N__7130),
            .I(N__7124));
    LocalMux I__948 (
            .O(N__7127),
            .I(N__7121));
    LocalMux I__947 (
            .O(N__7124),
            .I(\d1.countZ0Z_14 ));
    Odrv4 I__946 (
            .O(N__7121),
            .I(\d1.countZ0Z_14 ));
    InMux I__945 (
            .O(N__7116),
            .I(\d1.un3_count_cry_13 ));
    InMux I__944 (
            .O(N__7113),
            .I(N__7108));
    InMux I__943 (
            .O(N__7112),
            .I(N__7103));
    InMux I__942 (
            .O(N__7111),
            .I(N__7103));
    LocalMux I__941 (
            .O(N__7108),
            .I(\d1.countZ0Z_15 ));
    LocalMux I__940 (
            .O(N__7103),
            .I(\d1.countZ0Z_15 ));
    InMux I__939 (
            .O(N__7098),
            .I(\d1.un3_count_cry_14 ));
    InMux I__938 (
            .O(N__7095),
            .I(\d1.un3_count_cry_15 ));
    CascadeMux I__937 (
            .O(N__7092),
            .I(N__7087));
    InMux I__936 (
            .O(N__7091),
            .I(N__7084));
    InMux I__935 (
            .O(N__7090),
            .I(N__7079));
    InMux I__934 (
            .O(N__7087),
            .I(N__7079));
    LocalMux I__933 (
            .O(N__7084),
            .I(\d1.countZ0Z_16 ));
    LocalMux I__932 (
            .O(N__7079),
            .I(\d1.countZ0Z_16 ));
    SRMux I__931 (
            .O(N__7074),
            .I(N__7062));
    SRMux I__930 (
            .O(N__7073),
            .I(N__7062));
    SRMux I__929 (
            .O(N__7072),
            .I(N__7062));
    SRMux I__928 (
            .O(N__7071),
            .I(N__7062));
    GlobalMux I__927 (
            .O(N__7062),
            .I(N__7059));
    gio2CtrlBuf I__926 (
            .O(N__7059),
            .I(\d1.idle_i_g ));
    InMux I__925 (
            .O(N__7056),
            .I(N__7053));
    LocalMux I__924 (
            .O(N__7053),
            .I(N__7050));
    Span4Mux_v I__923 (
            .O(N__7050),
            .I(N__7047));
    Span4Mux_h I__922 (
            .O(N__7047),
            .I(N__7044));
    Odrv4 I__921 (
            .O(N__7044),
            .I(switch_dn_c));
    CascadeMux I__920 (
            .O(N__7041),
            .I(N__7037));
    InMux I__919 (
            .O(N__7040),
            .I(N__7033));
    InMux I__918 (
            .O(N__7037),
            .I(N__7030));
    InMux I__917 (
            .O(N__7036),
            .I(N__7027));
    LocalMux I__916 (
            .O(N__7033),
            .I(\a.countZ0Z_1 ));
    LocalMux I__915 (
            .O(N__7030),
            .I(\a.countZ0Z_1 ));
    LocalMux I__914 (
            .O(N__7027),
            .I(\a.countZ0Z_1 ));
    InMux I__913 (
            .O(N__7020),
            .I(N__7016));
    InMux I__912 (
            .O(N__7019),
            .I(N__7013));
    LocalMux I__911 (
            .O(N__7016),
            .I(\a.countZ0Z_2 ));
    LocalMux I__910 (
            .O(N__7013),
            .I(\a.countZ0Z_2 ));
    InMux I__909 (
            .O(N__7008),
            .I(\a.count_1_cry_1 ));
    InMux I__908 (
            .O(N__7005),
            .I(N__7001));
    InMux I__907 (
            .O(N__7004),
            .I(N__6998));
    LocalMux I__906 (
            .O(N__7001),
            .I(\a.countZ0Z_3 ));
    LocalMux I__905 (
            .O(N__6998),
            .I(\a.countZ0Z_3 ));
    InMux I__904 (
            .O(N__6993),
            .I(\a.count_1_cry_2 ));
    InMux I__903 (
            .O(N__6990),
            .I(\d1.un3_count_cry_4 ));
    InMux I__902 (
            .O(N__6987),
            .I(\d1.un3_count_cry_5 ));
    InMux I__901 (
            .O(N__6984),
            .I(\d1.un3_count_cry_6 ));
    InMux I__900 (
            .O(N__6981),
            .I(\d1.un3_count_cry_7 ));
    InMux I__899 (
            .O(N__6978),
            .I(bfn_7_17_0_));
    InMux I__898 (
            .O(N__6975),
            .I(\d1.un3_count_cry_9 ));
    InMux I__897 (
            .O(N__6972),
            .I(\d1.un3_count_cry_10 ));
    InMux I__896 (
            .O(N__6969),
            .I(\d1.un3_count_cry_11 ));
    InMux I__895 (
            .O(N__6966),
            .I(N__6962));
    InMux I__894 (
            .O(N__6965),
            .I(N__6959));
    LocalMux I__893 (
            .O(N__6962),
            .I(N__6956));
    LocalMux I__892 (
            .O(N__6959),
            .I(\d1.countZ0Z_13 ));
    Odrv4 I__891 (
            .O(N__6956),
            .I(\d1.countZ0Z_13 ));
    InMux I__890 (
            .O(N__6951),
            .I(\d1.un3_count_cry_12 ));
    CascadeMux I__889 (
            .O(N__6948),
            .I(N__6945));
    InMux I__888 (
            .O(N__6945),
            .I(N__6941));
    InMux I__887 (
            .O(N__6944),
            .I(N__6938));
    LocalMux I__886 (
            .O(N__6941),
            .I(N__6935));
    LocalMux I__885 (
            .O(N__6938),
            .I(\d1.syncZ0Z_1 ));
    Odrv4 I__884 (
            .O(N__6935),
            .I(\d1.syncZ0Z_1 ));
    CascadeMux I__883 (
            .O(N__6930),
            .I(\d1.trans_up_1_12_cascade_ ));
    InMux I__882 (
            .O(N__6927),
            .I(N__6924));
    LocalMux I__881 (
            .O(N__6924),
            .I(\d1.g1_3 ));
    CascadeMux I__880 (
            .O(N__6921),
            .I(\d1.g1_4_cascade_ ));
    CascadeMux I__879 (
            .O(N__6918),
            .I(N__6914));
    InMux I__878 (
            .O(N__6917),
            .I(N__6909));
    InMux I__877 (
            .O(N__6914),
            .I(N__6906));
    InMux I__876 (
            .O(N__6913),
            .I(N__6901));
    InMux I__875 (
            .O(N__6912),
            .I(N__6901));
    LocalMux I__874 (
            .O(N__6909),
            .I(\d1.countZ0Z_1 ));
    LocalMux I__873 (
            .O(N__6906),
            .I(\d1.countZ0Z_1 ));
    LocalMux I__872 (
            .O(N__6901),
            .I(\d1.countZ0Z_1 ));
    CascadeMux I__871 (
            .O(N__6894),
            .I(N__6890));
    InMux I__870 (
            .O(N__6893),
            .I(N__6886));
    InMux I__869 (
            .O(N__6890),
            .I(N__6881));
    InMux I__868 (
            .O(N__6889),
            .I(N__6881));
    LocalMux I__867 (
            .O(N__6886),
            .I(\d1.countZ0Z_2 ));
    LocalMux I__866 (
            .O(N__6881),
            .I(\d1.countZ0Z_2 ));
    InMux I__865 (
            .O(N__6876),
            .I(\d1.un3_count_cry_1 ));
    InMux I__864 (
            .O(N__6873),
            .I(\d1.un3_count_cry_2 ));
    InMux I__863 (
            .O(N__6870),
            .I(\d1.un3_count_cry_3 ));
    InMux I__862 (
            .O(N__6867),
            .I(N__6849));
    InMux I__861 (
            .O(N__6866),
            .I(N__6849));
    InMux I__860 (
            .O(N__6865),
            .I(N__6849));
    InMux I__859 (
            .O(N__6864),
            .I(N__6849));
    InMux I__858 (
            .O(N__6863),
            .I(N__6849));
    InMux I__857 (
            .O(N__6862),
            .I(N__6849));
    LocalMux I__856 (
            .O(N__6849),
            .I(\a.BUZZER3_20 ));
    CascadeMux I__855 (
            .O(N__6846),
            .I(N__6837));
    CascadeMux I__854 (
            .O(N__6845),
            .I(N__6834));
    CascadeMux I__853 (
            .O(N__6844),
            .I(N__6831));
    CascadeMux I__852 (
            .O(N__6843),
            .I(N__6828));
    CascadeMux I__851 (
            .O(N__6842),
            .I(N__6825));
    CascadeMux I__850 (
            .O(N__6841),
            .I(N__6822));
    InMux I__849 (
            .O(N__6840),
            .I(N__6819));
    InMux I__848 (
            .O(N__6837),
            .I(N__6810));
    InMux I__847 (
            .O(N__6834),
            .I(N__6810));
    InMux I__846 (
            .O(N__6831),
            .I(N__6810));
    InMux I__845 (
            .O(N__6828),
            .I(N__6810));
    InMux I__844 (
            .O(N__6825),
            .I(N__6805));
    InMux I__843 (
            .O(N__6822),
            .I(N__6805));
    LocalMux I__842 (
            .O(N__6819),
            .I(\a.BUZZER3_19 ));
    LocalMux I__841 (
            .O(N__6810),
            .I(\a.BUZZER3_19 ));
    LocalMux I__840 (
            .O(N__6805),
            .I(\a.BUZZER3_19 ));
    InMux I__839 (
            .O(N__6798),
            .I(N__6795));
    LocalMux I__838 (
            .O(N__6795),
            .I(\a.BUZZER3_18 ));
    InMux I__837 (
            .O(N__6792),
            .I(N__6789));
    LocalMux I__836 (
            .O(N__6789),
            .I(\a.BUZZER3_17 ));
    CascadeMux I__835 (
            .O(N__6786),
            .I(\a.BUZZER3_16_cascade_ ));
    InMux I__834 (
            .O(N__6783),
            .I(N__6780));
    LocalMux I__833 (
            .O(N__6780),
            .I(N__6771));
    InMux I__832 (
            .O(N__6779),
            .I(N__6758));
    InMux I__831 (
            .O(N__6778),
            .I(N__6758));
    InMux I__830 (
            .O(N__6777),
            .I(N__6758));
    InMux I__829 (
            .O(N__6776),
            .I(N__6758));
    InMux I__828 (
            .O(N__6775),
            .I(N__6758));
    InMux I__827 (
            .O(N__6774),
            .I(N__6758));
    Odrv4 I__826 (
            .O(N__6771),
            .I(\a.BUZZER3_24 ));
    LocalMux I__825 (
            .O(N__6758),
            .I(\a.BUZZER3_24 ));
    CascadeMux I__824 (
            .O(N__6753),
            .I(\a.BUZZER3_14_cascade_ ));
    CascadeMux I__823 (
            .O(N__6750),
            .I(\a.BUZZER3_20_cascade_ ));
    IoInMux I__822 (
            .O(N__6747),
            .I(N__6744));
    LocalMux I__821 (
            .O(N__6744),
            .I(N__6741));
    Span12Mux_s10_h I__820 (
            .O(N__6741),
            .I(N__6738));
    Span12Mux_v I__819 (
            .O(N__6738),
            .I(N__6734));
    InMux I__818 (
            .O(N__6737),
            .I(N__6731));
    Odrv12 I__817 (
            .O(N__6734),
            .I(BUZZER_c));
    LocalMux I__816 (
            .O(N__6731),
            .I(BUZZER_c));
    CascadeMux I__815 (
            .O(N__6726),
            .I(N__6723));
    InMux I__814 (
            .O(N__6723),
            .I(N__6719));
    InMux I__813 (
            .O(N__6722),
            .I(N__6716));
    LocalMux I__812 (
            .O(N__6719),
            .I(N__6713));
    LocalMux I__811 (
            .O(N__6716),
            .I(\display1.prescalerZ0Z_22 ));
    Odrv4 I__810 (
            .O(N__6713),
            .I(\display1.prescalerZ0Z_22 ));
    InMux I__809 (
            .O(N__6708),
            .I(\display1.prescaler_2_cry_21 ));
    InMux I__808 (
            .O(N__6705),
            .I(\display1.prescaler_2_cry_22 ));
    CascadeMux I__807 (
            .O(N__6702),
            .I(N__6699));
    InMux I__806 (
            .O(N__6699),
            .I(N__6696));
    LocalMux I__805 (
            .O(N__6696),
            .I(N__6692));
    InMux I__804 (
            .O(N__6695),
            .I(N__6689));
    Span4Mux_h I__803 (
            .O(N__6692),
            .I(N__6686));
    LocalMux I__802 (
            .O(N__6689),
            .I(\display1.prescalerZ0Z_23 ));
    Odrv4 I__801 (
            .O(N__6686),
            .I(\display1.prescalerZ0Z_23 ));
    InMux I__800 (
            .O(N__6681),
            .I(N__6677));
    InMux I__799 (
            .O(N__6680),
            .I(N__6674));
    LocalMux I__798 (
            .O(N__6677),
            .I(\display1.prescalerZ0Z_12 ));
    LocalMux I__797 (
            .O(N__6674),
            .I(\display1.prescalerZ0Z_12 ));
    InMux I__796 (
            .O(N__6669),
            .I(N__6665));
    InMux I__795 (
            .O(N__6668),
            .I(N__6662));
    LocalMux I__794 (
            .O(N__6665),
            .I(\display1.prescalerZ0Z_11 ));
    LocalMux I__793 (
            .O(N__6662),
            .I(\display1.prescalerZ0Z_11 ));
    CascadeMux I__792 (
            .O(N__6657),
            .I(N__6653));
    InMux I__791 (
            .O(N__6656),
            .I(N__6650));
    InMux I__790 (
            .O(N__6653),
            .I(N__6647));
    LocalMux I__789 (
            .O(N__6650),
            .I(\display1.prescalerZ0Z_13 ));
    LocalMux I__788 (
            .O(N__6647),
            .I(\display1.prescalerZ0Z_13 ));
    InMux I__787 (
            .O(N__6642),
            .I(N__6638));
    InMux I__786 (
            .O(N__6641),
            .I(N__6635));
    LocalMux I__785 (
            .O(N__6638),
            .I(\display1.prescalerZ0Z_10 ));
    LocalMux I__784 (
            .O(N__6635),
            .I(\display1.prescalerZ0Z_10 ));
    InMux I__783 (
            .O(N__6630),
            .I(N__6627));
    LocalMux I__782 (
            .O(N__6627),
            .I(N__6624));
    Span4Mux_h I__781 (
            .O(N__6624),
            .I(N__6621));
    Odrv4 I__780 (
            .O(N__6621),
            .I(\display1.prescaler8_12 ));
    IoInMux I__779 (
            .O(N__6618),
            .I(N__6615));
    LocalMux I__778 (
            .O(N__6615),
            .I(N__6612));
    Span12Mux_s9_h I__777 (
            .O(N__6612),
            .I(N__6609));
    Odrv12 I__776 (
            .O(N__6609),
            .I(\d1.idle_i ));
    CascadeMux I__775 (
            .O(N__6606),
            .I(\d1.trans_up_1_11_cascade_ ));
    InMux I__774 (
            .O(N__6603),
            .I(N__6600));
    LocalMux I__773 (
            .O(N__6600),
            .I(N__6596));
    InMux I__772 (
            .O(N__6599),
            .I(N__6593));
    Odrv4 I__771 (
            .O(N__6596),
            .I(\display1.prescalerZ0Z_14 ));
    LocalMux I__770 (
            .O(N__6593),
            .I(\display1.prescalerZ0Z_14 ));
    InMux I__769 (
            .O(N__6588),
            .I(N__6585));
    LocalMux I__768 (
            .O(N__6585),
            .I(N__6582));
    Odrv4 I__767 (
            .O(N__6582),
            .I(\display1.prescaler_2_14 ));
    InMux I__766 (
            .O(N__6579),
            .I(\display1.prescaler_2_cry_13 ));
    CascadeMux I__765 (
            .O(N__6576),
            .I(N__6572));
    InMux I__764 (
            .O(N__6575),
            .I(N__6569));
    InMux I__763 (
            .O(N__6572),
            .I(N__6566));
    LocalMux I__762 (
            .O(N__6569),
            .I(N__6563));
    LocalMux I__761 (
            .O(N__6566),
            .I(N__6560));
    Odrv12 I__760 (
            .O(N__6563),
            .I(\display1.prescalerZ0Z_15 ));
    Odrv4 I__759 (
            .O(N__6560),
            .I(\display1.prescalerZ0Z_15 ));
    InMux I__758 (
            .O(N__6555),
            .I(N__6552));
    LocalMux I__757 (
            .O(N__6552),
            .I(N__6549));
    Odrv4 I__756 (
            .O(N__6549),
            .I(\display1.prescaler_2_15 ));
    InMux I__755 (
            .O(N__6546),
            .I(\display1.prescaler_2_cry_14 ));
    InMux I__754 (
            .O(N__6543),
            .I(N__6539));
    InMux I__753 (
            .O(N__6542),
            .I(N__6536));
    LocalMux I__752 (
            .O(N__6539),
            .I(N__6533));
    LocalMux I__751 (
            .O(N__6536),
            .I(\display1.prescalerZ0Z_16 ));
    Odrv4 I__750 (
            .O(N__6533),
            .I(\display1.prescalerZ0Z_16 ));
    InMux I__749 (
            .O(N__6528),
            .I(\display1.prescaler_2_cry_15 ));
    InMux I__748 (
            .O(N__6525),
            .I(N__6521));
    InMux I__747 (
            .O(N__6524),
            .I(N__6518));
    LocalMux I__746 (
            .O(N__6521),
            .I(N__6515));
    LocalMux I__745 (
            .O(N__6518),
            .I(N__6510));
    Span4Mux_v I__744 (
            .O(N__6515),
            .I(N__6510));
    Odrv4 I__743 (
            .O(N__6510),
            .I(\display1.prescalerZ0Z_17 ));
    InMux I__742 (
            .O(N__6507),
            .I(bfn_5_15_0_));
    CascadeMux I__741 (
            .O(N__6504),
            .I(N__6501));
    InMux I__740 (
            .O(N__6501),
            .I(N__6498));
    LocalMux I__739 (
            .O(N__6498),
            .I(N__6494));
    InMux I__738 (
            .O(N__6497),
            .I(N__6491));
    Span4Mux_v I__737 (
            .O(N__6494),
            .I(N__6488));
    LocalMux I__736 (
            .O(N__6491),
            .I(\display1.prescalerZ0Z_18 ));
    Odrv4 I__735 (
            .O(N__6488),
            .I(\display1.prescalerZ0Z_18 ));
    InMux I__734 (
            .O(N__6483),
            .I(\display1.prescaler_2_cry_17 ));
    InMux I__733 (
            .O(N__6480),
            .I(N__6476));
    InMux I__732 (
            .O(N__6479),
            .I(N__6473));
    LocalMux I__731 (
            .O(N__6476),
            .I(N__6470));
    LocalMux I__730 (
            .O(N__6473),
            .I(\display1.prescalerZ0Z_19 ));
    Odrv4 I__729 (
            .O(N__6470),
            .I(\display1.prescalerZ0Z_19 ));
    InMux I__728 (
            .O(N__6465),
            .I(\display1.prescaler_2_cry_18 ));
    InMux I__727 (
            .O(N__6462),
            .I(N__6458));
    InMux I__726 (
            .O(N__6461),
            .I(N__6455));
    LocalMux I__725 (
            .O(N__6458),
            .I(N__6452));
    LocalMux I__724 (
            .O(N__6455),
            .I(\display1.prescalerZ0Z_20 ));
    Odrv4 I__723 (
            .O(N__6452),
            .I(\display1.prescalerZ0Z_20 ));
    InMux I__722 (
            .O(N__6447),
            .I(\display1.prescaler_2_cry_19 ));
    InMux I__721 (
            .O(N__6444),
            .I(N__6440));
    InMux I__720 (
            .O(N__6443),
            .I(N__6437));
    LocalMux I__719 (
            .O(N__6440),
            .I(N__6434));
    LocalMux I__718 (
            .O(N__6437),
            .I(\display1.prescalerZ0Z_21 ));
    Odrv4 I__717 (
            .O(N__6434),
            .I(\display1.prescalerZ0Z_21 ));
    InMux I__716 (
            .O(N__6429),
            .I(\display1.prescaler_2_cry_20 ));
    InMux I__715 (
            .O(N__6426),
            .I(N__6423));
    LocalMux I__714 (
            .O(N__6423),
            .I(N__6419));
    InMux I__713 (
            .O(N__6422),
            .I(N__6416));
    Odrv4 I__712 (
            .O(N__6419),
            .I(\display1.prescalerZ0Z_6 ));
    LocalMux I__711 (
            .O(N__6416),
            .I(\display1.prescalerZ0Z_6 ));
    InMux I__710 (
            .O(N__6411),
            .I(N__6408));
    LocalMux I__709 (
            .O(N__6408),
            .I(N__6405));
    Odrv4 I__708 (
            .O(N__6405),
            .I(\display1.prescaler_2_6 ));
    InMux I__707 (
            .O(N__6402),
            .I(\display1.prescaler_2_cry_5 ));
    CascadeMux I__706 (
            .O(N__6399),
            .I(N__6395));
    InMux I__705 (
            .O(N__6398),
            .I(N__6392));
    InMux I__704 (
            .O(N__6395),
            .I(N__6389));
    LocalMux I__703 (
            .O(N__6392),
            .I(\display1.prescalerZ0Z_7 ));
    LocalMux I__702 (
            .O(N__6389),
            .I(\display1.prescalerZ0Z_7 ));
    InMux I__701 (
            .O(N__6384),
            .I(\display1.prescaler_2_cry_6 ));
    InMux I__700 (
            .O(N__6381),
            .I(N__6378));
    LocalMux I__699 (
            .O(N__6378),
            .I(N__6374));
    InMux I__698 (
            .O(N__6377),
            .I(N__6371));
    Odrv4 I__697 (
            .O(N__6374),
            .I(\display1.prescalerZ0Z_8 ));
    LocalMux I__696 (
            .O(N__6371),
            .I(\display1.prescalerZ0Z_8 ));
    InMux I__695 (
            .O(N__6366),
            .I(N__6363));
    LocalMux I__694 (
            .O(N__6363),
            .I(N__6360));
    Odrv4 I__693 (
            .O(N__6360),
            .I(\display1.prescaler_2_8 ));
    InMux I__692 (
            .O(N__6357),
            .I(\display1.prescaler_2_cry_7 ));
    InMux I__691 (
            .O(N__6354),
            .I(N__6351));
    LocalMux I__690 (
            .O(N__6351),
            .I(N__6347));
    InMux I__689 (
            .O(N__6350),
            .I(N__6344));
    Odrv4 I__688 (
            .O(N__6347),
            .I(\display1.prescalerZ0Z_9 ));
    LocalMux I__687 (
            .O(N__6344),
            .I(\display1.prescalerZ0Z_9 ));
    InMux I__686 (
            .O(N__6339),
            .I(N__6336));
    LocalMux I__685 (
            .O(N__6336),
            .I(N__6333));
    Odrv4 I__684 (
            .O(N__6333),
            .I(\display1.prescaler_2_9 ));
    InMux I__683 (
            .O(N__6330),
            .I(bfn_5_14_0_));
    InMux I__682 (
            .O(N__6327),
            .I(\display1.prescaler_2_cry_9 ));
    InMux I__681 (
            .O(N__6324),
            .I(\display1.prescaler_2_cry_10 ));
    InMux I__680 (
            .O(N__6321),
            .I(\display1.prescaler_2_cry_11 ));
    InMux I__679 (
            .O(N__6318),
            .I(\display1.prescaler_2_cry_12 ));
    CascadeMux I__678 (
            .O(N__6315),
            .I(\display1.prescaler8_17_cascade_ ));
    InMux I__677 (
            .O(N__6312),
            .I(N__6298));
    InMux I__676 (
            .O(N__6311),
            .I(N__6298));
    InMux I__675 (
            .O(N__6310),
            .I(N__6298));
    InMux I__674 (
            .O(N__6309),
            .I(N__6291));
    InMux I__673 (
            .O(N__6308),
            .I(N__6291));
    InMux I__672 (
            .O(N__6307),
            .I(N__6291));
    InMux I__671 (
            .O(N__6306),
            .I(N__6286));
    InMux I__670 (
            .O(N__6305),
            .I(N__6286));
    LocalMux I__669 (
            .O(N__6298),
            .I(\display1.prescaler8_21 ));
    LocalMux I__668 (
            .O(N__6291),
            .I(\display1.prescaler8_21 ));
    LocalMux I__667 (
            .O(N__6286),
            .I(\display1.prescaler8_21 ));
    CascadeMux I__666 (
            .O(N__6279),
            .I(N__6274));
    CascadeMux I__665 (
            .O(N__6278),
            .I(N__6268));
    CascadeMux I__664 (
            .O(N__6277),
            .I(N__6265));
    InMux I__663 (
            .O(N__6274),
            .I(N__6256));
    InMux I__662 (
            .O(N__6273),
            .I(N__6256));
    InMux I__661 (
            .O(N__6272),
            .I(N__6256));
    InMux I__660 (
            .O(N__6271),
            .I(N__6256));
    InMux I__659 (
            .O(N__6268),
            .I(N__6249));
    InMux I__658 (
            .O(N__6265),
            .I(N__6249));
    LocalMux I__657 (
            .O(N__6256),
            .I(N__6246));
    InMux I__656 (
            .O(N__6255),
            .I(N__6241));
    InMux I__655 (
            .O(N__6254),
            .I(N__6241));
    LocalMux I__654 (
            .O(N__6249),
            .I(\display1.prescaler8_17 ));
    Odrv4 I__653 (
            .O(N__6246),
            .I(\display1.prescaler8_17 ));
    LocalMux I__652 (
            .O(N__6241),
            .I(\display1.prescaler8_17 ));
    CascadeMux I__651 (
            .O(N__6234),
            .I(N__6230));
    CascadeMux I__650 (
            .O(N__6233),
            .I(N__6227));
    InMux I__649 (
            .O(N__6230),
            .I(N__6215));
    InMux I__648 (
            .O(N__6227),
            .I(N__6215));
    InMux I__647 (
            .O(N__6226),
            .I(N__6215));
    InMux I__646 (
            .O(N__6225),
            .I(N__6212));
    InMux I__645 (
            .O(N__6224),
            .I(N__6205));
    InMux I__644 (
            .O(N__6223),
            .I(N__6205));
    InMux I__643 (
            .O(N__6222),
            .I(N__6205));
    LocalMux I__642 (
            .O(N__6215),
            .I(N__6198));
    LocalMux I__641 (
            .O(N__6212),
            .I(N__6198));
    LocalMux I__640 (
            .O(N__6205),
            .I(N__6195));
    InMux I__639 (
            .O(N__6204),
            .I(N__6190));
    InMux I__638 (
            .O(N__6203),
            .I(N__6190));
    Odrv4 I__637 (
            .O(N__6198),
            .I(\display1.prescaler8_16 ));
    Odrv4 I__636 (
            .O(N__6195),
            .I(\display1.prescaler8_16 ));
    LocalMux I__635 (
            .O(N__6190),
            .I(\display1.prescaler8_16 ));
    InMux I__634 (
            .O(N__6183),
            .I(N__6180));
    LocalMux I__633 (
            .O(N__6180),
            .I(N__6177));
    Span4Mux_h I__632 (
            .O(N__6177),
            .I(N__6174));
    Odrv4 I__631 (
            .O(N__6174),
            .I(\display1.prescaler8_13 ));
    InMux I__630 (
            .O(N__6171),
            .I(N__6168));
    LocalMux I__629 (
            .O(N__6168),
            .I(N__6163));
    InMux I__628 (
            .O(N__6167),
            .I(N__6158));
    InMux I__627 (
            .O(N__6166),
            .I(N__6158));
    Odrv4 I__626 (
            .O(N__6163),
            .I(\display1.prescalerZ0Z_1 ));
    LocalMux I__625 (
            .O(N__6158),
            .I(\display1.prescalerZ0Z_1 ));
    CascadeMux I__624 (
            .O(N__6153),
            .I(N__6150));
    InMux I__623 (
            .O(N__6150),
            .I(N__6144));
    InMux I__622 (
            .O(N__6149),
            .I(N__6139));
    InMux I__621 (
            .O(N__6148),
            .I(N__6139));
    InMux I__620 (
            .O(N__6147),
            .I(N__6136));
    LocalMux I__619 (
            .O(N__6144),
            .I(N__6133));
    LocalMux I__618 (
            .O(N__6139),
            .I(\display1.prescalerZ0Z_0 ));
    LocalMux I__617 (
            .O(N__6136),
            .I(\display1.prescalerZ0Z_0 ));
    Odrv12 I__616 (
            .O(N__6133),
            .I(\display1.prescalerZ0Z_0 ));
    InMux I__615 (
            .O(N__6126),
            .I(N__6122));
    InMux I__614 (
            .O(N__6125),
            .I(N__6119));
    LocalMux I__613 (
            .O(N__6122),
            .I(\display1.prescalerZ0Z_2 ));
    LocalMux I__612 (
            .O(N__6119),
            .I(\display1.prescalerZ0Z_2 ));
    InMux I__611 (
            .O(N__6114),
            .I(\display1.prescaler_2_cry_1 ));
    InMux I__610 (
            .O(N__6111),
            .I(N__6107));
    InMux I__609 (
            .O(N__6110),
            .I(N__6104));
    LocalMux I__608 (
            .O(N__6107),
            .I(\display1.prescalerZ0Z_3 ));
    LocalMux I__607 (
            .O(N__6104),
            .I(\display1.prescalerZ0Z_3 ));
    InMux I__606 (
            .O(N__6099),
            .I(\display1.prescaler_2_cry_2 ));
    InMux I__605 (
            .O(N__6096),
            .I(N__6093));
    LocalMux I__604 (
            .O(N__6093),
            .I(N__6089));
    InMux I__603 (
            .O(N__6092),
            .I(N__6086));
    Odrv4 I__602 (
            .O(N__6089),
            .I(\display1.prescalerZ0Z_4 ));
    LocalMux I__601 (
            .O(N__6086),
            .I(\display1.prescalerZ0Z_4 ));
    InMux I__600 (
            .O(N__6081),
            .I(N__6078));
    LocalMux I__599 (
            .O(N__6078),
            .I(N__6075));
    Span4Mux_h I__598 (
            .O(N__6075),
            .I(N__6072));
    Odrv4 I__597 (
            .O(N__6072),
            .I(\display1.prescaler_2_4 ));
    InMux I__596 (
            .O(N__6069),
            .I(\display1.prescaler_2_cry_3 ));
    InMux I__595 (
            .O(N__6066),
            .I(N__6062));
    InMux I__594 (
            .O(N__6065),
            .I(N__6059));
    LocalMux I__593 (
            .O(N__6062),
            .I(\display1.prescalerZ0Z_5 ));
    LocalMux I__592 (
            .O(N__6059),
            .I(\display1.prescalerZ0Z_5 ));
    InMux I__591 (
            .O(N__6054),
            .I(\display1.prescaler_2_cry_4 ));
    InMux I__590 (
            .O(N__6051),
            .I(N__6048));
    LocalMux I__589 (
            .O(N__6048),
            .I(\display1.prescaler8_14 ));
    CascadeMux I__588 (
            .O(N__6045),
            .I(\display1.prescaler8_15_cascade_ ));
    CascadeMux I__587 (
            .O(N__6042),
            .I(\display1.prescaler8_21_cascade_ ));
    IoInMux I__586 (
            .O(N__6039),
            .I(N__6036));
    LocalMux I__585 (
            .O(N__6036),
            .I(N__6033));
    Span12Mux_s4_h I__584 (
            .O(N__6033),
            .I(N__6030));
    Odrv12 I__583 (
            .O(N__6030),
            .I(SEG1_c_2));
    IoInMux I__582 (
            .O(N__6027),
            .I(N__6024));
    LocalMux I__581 (
            .O(N__6024),
            .I(N__6021));
    IoSpan4Mux I__580 (
            .O(N__6021),
            .I(N__6018));
    Span4Mux_s3_v I__579 (
            .O(N__6018),
            .I(N__6015));
    Span4Mux_v I__578 (
            .O(N__6015),
            .I(N__6012));
    Span4Mux_v I__577 (
            .O(N__6012),
            .I(N__6009));
    Odrv4 I__576 (
            .O(N__6009),
            .I(SEG1_c_0));
    CascadeMux I__575 (
            .O(N__6006),
            .I(\display1.prescaler8_cascade_ ));
    CascadeMux I__574 (
            .O(N__6003),
            .I(N__5997));
    CascadeMux I__573 (
            .O(N__6002),
            .I(N__5994));
    CascadeMux I__572 (
            .O(N__6001),
            .I(N__5990));
    CascadeMux I__571 (
            .O(N__6000),
            .I(N__5987));
    InMux I__570 (
            .O(N__5997),
            .I(N__5977));
    InMux I__569 (
            .O(N__5994),
            .I(N__5977));
    InMux I__568 (
            .O(N__5993),
            .I(N__5977));
    InMux I__567 (
            .O(N__5990),
            .I(N__5968));
    InMux I__566 (
            .O(N__5987),
            .I(N__5968));
    InMux I__565 (
            .O(N__5986),
            .I(N__5968));
    InMux I__564 (
            .O(N__5985),
            .I(N__5968));
    InMux I__563 (
            .O(N__5984),
            .I(N__5965));
    LocalMux I__562 (
            .O(N__5977),
            .I(\display1.digit_dataZ0Z_3 ));
    LocalMux I__561 (
            .O(N__5968),
            .I(\display1.digit_dataZ0Z_3 ));
    LocalMux I__560 (
            .O(N__5965),
            .I(\display1.digit_dataZ0Z_3 ));
    IoInMux I__559 (
            .O(N__5958),
            .I(N__5955));
    LocalMux I__558 (
            .O(N__5955),
            .I(N__5952));
    IoSpan4Mux I__557 (
            .O(N__5952),
            .I(N__5949));
    Span4Mux_s3_h I__556 (
            .O(N__5949),
            .I(N__5946));
    Span4Mux_v I__555 (
            .O(N__5946),
            .I(N__5943));
    Span4Mux_v I__554 (
            .O(N__5943),
            .I(N__5940));
    Odrv4 I__553 (
            .O(N__5940),
            .I(DIGIT_c_0));
    CascadeMux I__552 (
            .O(N__5937),
            .I(N__5932));
    CascadeMux I__551 (
            .O(N__5936),
            .I(N__5927));
    CascadeMux I__550 (
            .O(N__5935),
            .I(N__5922));
    InMux I__549 (
            .O(N__5932),
            .I(N__5913));
    InMux I__548 (
            .O(N__5931),
            .I(N__5913));
    InMux I__547 (
            .O(N__5930),
            .I(N__5913));
    InMux I__546 (
            .O(N__5927),
            .I(N__5913));
    InMux I__545 (
            .O(N__5926),
            .I(N__5906));
    InMux I__544 (
            .O(N__5925),
            .I(N__5906));
    InMux I__543 (
            .O(N__5922),
            .I(N__5906));
    LocalMux I__542 (
            .O(N__5913),
            .I(\display1.digit_dataZ0Z_2 ));
    LocalMux I__541 (
            .O(N__5906),
            .I(\display1.digit_dataZ0Z_2 ));
    InMux I__540 (
            .O(N__5901),
            .I(N__5886));
    InMux I__539 (
            .O(N__5900),
            .I(N__5886));
    InMux I__538 (
            .O(N__5899),
            .I(N__5886));
    InMux I__537 (
            .O(N__5898),
            .I(N__5886));
    InMux I__536 (
            .O(N__5897),
            .I(N__5879));
    InMux I__535 (
            .O(N__5896),
            .I(N__5879));
    InMux I__534 (
            .O(N__5895),
            .I(N__5879));
    LocalMux I__533 (
            .O(N__5886),
            .I(\display1.digit_dataZ0Z_1 ));
    LocalMux I__532 (
            .O(N__5879),
            .I(\display1.digit_dataZ0Z_1 ));
    CascadeMux I__531 (
            .O(N__5874),
            .I(N__5866));
    InMux I__530 (
            .O(N__5873),
            .I(N__5863));
    InMux I__529 (
            .O(N__5872),
            .I(N__5854));
    InMux I__528 (
            .O(N__5871),
            .I(N__5854));
    InMux I__527 (
            .O(N__5870),
            .I(N__5854));
    InMux I__526 (
            .O(N__5869),
            .I(N__5854));
    InMux I__525 (
            .O(N__5866),
            .I(N__5851));
    LocalMux I__524 (
            .O(N__5863),
            .I(\display1.digit_posnZ0 ));
    LocalMux I__523 (
            .O(N__5854),
            .I(\display1.digit_posnZ0 ));
    LocalMux I__522 (
            .O(N__5851),
            .I(\display1.digit_posnZ0 ));
    InMux I__521 (
            .O(N__5844),
            .I(N__5829));
    InMux I__520 (
            .O(N__5843),
            .I(N__5829));
    InMux I__519 (
            .O(N__5842),
            .I(N__5829));
    InMux I__518 (
            .O(N__5841),
            .I(N__5829));
    InMux I__517 (
            .O(N__5840),
            .I(N__5822));
    InMux I__516 (
            .O(N__5839),
            .I(N__5822));
    InMux I__515 (
            .O(N__5838),
            .I(N__5822));
    LocalMux I__514 (
            .O(N__5829),
            .I(\display1.digit_dataZ0Z_0 ));
    LocalMux I__513 (
            .O(N__5822),
            .I(\display1.digit_dataZ0Z_0 ));
    CEMux I__512 (
            .O(N__5817),
            .I(N__5814));
    LocalMux I__511 (
            .O(N__5814),
            .I(\display1.prescaler8 ));
    IoInMux I__510 (
            .O(N__5811),
            .I(N__5808));
    LocalMux I__509 (
            .O(N__5808),
            .I(N__5805));
    IoSpan4Mux I__508 (
            .O(N__5805),
            .I(N__5802));
    Span4Mux_s1_h I__507 (
            .O(N__5802),
            .I(N__5799));
    Odrv4 I__506 (
            .O(N__5799),
            .I(SEG1_c_5));
    IoInMux I__505 (
            .O(N__5796),
            .I(N__5793));
    LocalMux I__504 (
            .O(N__5793),
            .I(N__5790));
    IoSpan4Mux I__503 (
            .O(N__5790),
            .I(N__5787));
    Span4Mux_s3_h I__502 (
            .O(N__5787),
            .I(N__5784));
    Odrv4 I__501 (
            .O(N__5784),
            .I(SEG1_c_6));
    IoInMux I__500 (
            .O(N__5781),
            .I(N__5778));
    LocalMux I__499 (
            .O(N__5778),
            .I(N__5775));
    Odrv12 I__498 (
            .O(N__5775),
            .I(SEG1_c_4));
    IoInMux I__497 (
            .O(N__5772),
            .I(N__5769));
    LocalMux I__496 (
            .O(N__5769),
            .I(N__5766));
    Odrv12 I__495 (
            .O(N__5766),
            .I(SEG1_c_3));
    IoInMux I__494 (
            .O(N__5763),
            .I(N__5760));
    LocalMux I__493 (
            .O(N__5760),
            .I(N__5757));
    Span4Mux_s3_h I__492 (
            .O(N__5757),
            .I(N__5754));
    Span4Mux_v I__491 (
            .O(N__5754),
            .I(N__5751));
    Odrv4 I__490 (
            .O(N__5751),
            .I(SEG1_c_1));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(prescaler_1_cry_8),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(prescaler_1_cry_16),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(prescaler_1_cry_24),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\display2.prescaler_2_cry_8 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\display2.prescaler_2_cry_16 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\display1.prescaler_2_cry_8 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\display1.prescaler_2_cry_16 ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\d4.un3_count_cry_8 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\d3.un3_count_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\d2.un3_count_cry_8 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(\d1.un3_count_cry_8 ),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\a.count_1_cry_8 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\a.count_1_cry_16 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\a.count_1_cry_24 ),
            .carryinitout(bfn_8_14_0_));
    ICE_GB un1_state_3_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__10560),
            .GLOBALBUFFEROUTPUT(un1_state_3_g));
    ICE_GB \d4.sync_1_RNIQPEK_0  (
            .USERSIGNALTOGLOBALBUFFER(N__8529),
            .GLOBALBUFFEROUTPUT(\d4.idle_i_g ));
    ICE_GB \d3.state_RNIOCAC_0  (
            .USERSIGNALTOGLOBALBUFFER(N__12543),
            .GLOBALBUFFEROUTPUT(\d3.idle_i_g ));
    ICE_GB \d2.sync_1_RNIMV5K_0  (
            .USERSIGNALTOGLOBALBUFFER(N__11928),
            .GLOBALBUFFEROUTPUT(\d2.idle_i_g ));
    ICE_GB \d1.sync_1_RNIKI1C_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6618),
            .GLOBALBUFFEROUTPUT(\d1.idle_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \display1.decoder.SEG_5_LC_1_14_2 .C_ON=1'b0;
    defparam \display1.decoder.SEG_5_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_5_LC_1_14_2 .LUT_INIT=16'b0000100100111111;
    LogicCell40 \display1.decoder.SEG_5_LC_1_14_2  (
            .in0(N__5843),
            .in1(N__5900),
            .in2(N__6001),
            .in3(N__5931),
            .lcout(SEG1_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14273),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_6_LC_1_14_3 .C_ON=1'b0;
    defparam \display1.decoder.SEG_6_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_6_LC_1_14_3 .LUT_INIT=16'b0011011000100111;
    LogicCell40 \display1.decoder.SEG_6_LC_1_14_3  (
            .in0(N__5901),
            .in1(N__5986),
            .in2(N__5937),
            .in3(N__5844),
            .lcout(SEG1_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14273),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_4_LC_1_14_4 .C_ON=1'b0;
    defparam \display1.decoder.SEG_4_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_4_LC_1_14_4 .LUT_INIT=16'b0000111100111011;
    LogicCell40 \display1.decoder.SEG_4_LC_1_14_4  (
            .in0(N__5842),
            .in1(N__5899),
            .in2(N__6000),
            .in3(N__5930),
            .lcout(SEG1_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14273),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_3_LC_1_14_7 .C_ON=1'b0;
    defparam \display1.decoder.SEG_3_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_3_LC_1_14_7 .LUT_INIT=16'b0001011000100111;
    LogicCell40 \display1.decoder.SEG_3_LC_1_14_7  (
            .in0(N__5898),
            .in1(N__5985),
            .in2(N__5936),
            .in3(N__5841),
            .lcout(SEG1_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14273),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_1_LC_1_15_0 .C_ON=1'b0;
    defparam \display1.decoder.SEG_1_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_1_LC_1_15_0 .LUT_INIT=16'b0000011100110001;
    LogicCell40 \display1.decoder.SEG_1_LC_1_15_0  (
            .in0(N__5839),
            .in1(N__5896),
            .in2(N__6002),
            .in3(N__5925),
            .lcout(SEG1_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14268),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_2_LC_1_15_4 .C_ON=1'b0;
    defparam \display1.decoder.SEG_2_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_2_LC_1_15_4 .LUT_INIT=16'b0000010000010101;
    LogicCell40 \display1.decoder.SEG_2_LC_1_15_4  (
            .in0(N__5840),
            .in1(N__5897),
            .in2(N__6003),
            .in3(N__5926),
            .lcout(SEG1_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14268),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.decoder.SEG_0_LC_1_15_7 .C_ON=1'b0;
    defparam \display1.decoder.SEG_0_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \display1.decoder.SEG_0_LC_1_15_7 .LUT_INIT=16'b0001011000110110;
    LogicCell40 \display1.decoder.SEG_0_LC_1_15_7  (
            .in0(N__5895),
            .in1(N__5993),
            .in2(N__5935),
            .in3(N__5838),
            .lcout(SEG1_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14268),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNI2HUD5_16_LC_2_14_2 .C_ON=1'b0;
    defparam \display1.prescaler_RNI2HUD5_16_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNI2HUD5_16_LC_2_14_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \display1.prescaler_RNI2HUD5_16_LC_2_14_2  (
            .in0(N__6254),
            .in1(N__6203),
            .in2(_gnd_net_),
            .in3(N__6305),
            .lcout(\display1.prescaler8 ),
            .ltout(\display1.prescaler8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.digit_data_3_LC_2_14_3 .C_ON=1'b0;
    defparam \display1.digit_data_3_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \display1.digit_data_3_LC_2_14_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \display1.digit_data_3_LC_2_14_3  (
            .in0(N__5873),
            .in1(N__5984),
            .in2(N__6006),
            .in3(N__10407),
            .lcout(\display1.digit_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14269),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.digit_posn_LC_2_14_6 .C_ON=1'b0;
    defparam \display1.digit_posn_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \display1.digit_posn_LC_2_14_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \display1.digit_posn_LC_2_14_6  (
            .in0(N__6255),
            .in1(N__6204),
            .in2(N__5874),
            .in3(N__6306),
            .lcout(\display1.digit_posnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14269),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.DIGIT_e_0_LC_2_15_4 .C_ON=1'b0;
    defparam \display1.DIGIT_e_0_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \display1.DIGIT_e_0_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \display1.DIGIT_e_0_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5872),
            .lcout(DIGIT_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14265),
            .ce(N__5817),
            .sr(_gnd_net_));
    defparam \display1.digit_data_e_0_2_LC_2_15_5 .C_ON=1'b0;
    defparam \display1.digit_data_e_0_2_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \display1.digit_data_e_0_2_LC_2_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \display1.digit_data_e_0_2_LC_2_15_5  (
            .in0(N__5871),
            .in1(N__10482),
            .in2(_gnd_net_),
            .in3(N__10600),
            .lcout(\display1.digit_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14265),
            .ce(N__5817),
            .sr(_gnd_net_));
    defparam \display1.digit_data_e_0_1_LC_2_15_6 .C_ON=1'b0;
    defparam \display1.digit_data_e_0_1_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \display1.digit_data_e_0_1_LC_2_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \display1.digit_data_e_0_1_LC_2_15_6  (
            .in0(N__10446),
            .in1(N__12507),
            .in2(_gnd_net_),
            .in3(N__5870),
            .lcout(\display1.digit_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14265),
            .ce(N__5817),
            .sr(_gnd_net_));
    defparam \display1.digit_data_e_0_0_LC_2_15_7 .C_ON=1'b0;
    defparam \display1.digit_data_e_0_0_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \display1.digit_data_e_0_0_LC_2_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \display1.digit_data_e_0_0_LC_2_15_7  (
            .in0(N__5869),
            .in1(N__10368),
            .in2(_gnd_net_),
            .in3(N__12456),
            .lcout(\display1.digit_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14265),
            .ce(N__5817),
            .sr(_gnd_net_));
    defparam \display1.prescaler_8_LC_3_13_0 .C_ON=1'b0;
    defparam \display1.prescaler_8_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_8_LC_3_13_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display1.prescaler_8_LC_3_13_0  (
            .in0(N__6309),
            .in1(N__6273),
            .in2(N__6234),
            .in3(N__6366),
            .lcout(\display1.prescalerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14270),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_4_LC_3_13_1 .C_ON=1'b0;
    defparam \display1.prescaler_4_LC_3_13_1 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_4_LC_3_13_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \display1.prescaler_4_LC_3_13_1  (
            .in0(N__6225),
            .in1(N__6081),
            .in2(N__6279),
            .in3(N__6307),
            .lcout(\display1.prescalerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14270),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNID8UQ_1_LC_3_13_2 .C_ON=1'b0;
    defparam \display1.prescaler_RNID8UQ_1_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNID8UQ_1_LC_3_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \display1.prescaler_RNID8UQ_1_LC_3_13_2  (
            .in0(N__6599),
            .in1(N__6350),
            .in2(N__6576),
            .in3(N__6166),
            .lcout(\display1.prescaler8_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNIVNSK_23_LC_3_13_3 .C_ON=1'b0;
    defparam \display1.prescaler_RNIVNSK_23_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNIVNSK_23_LC_3_13_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \display1.prescaler_RNIVNSK_23_LC_3_13_3  (
            .in0(N__6377),
            .in1(N__6422),
            .in2(N__6702),
            .in3(N__6092),
            .lcout(),
            .ltout(\display1.prescaler8_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNIN1N53_1_LC_3_13_4 .C_ON=1'b0;
    defparam \display1.prescaler_RNIN1N53_1_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNIN1N53_1_LC_3_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \display1.prescaler_RNIN1N53_1_LC_3_13_4  (
            .in0(N__6051),
            .in1(N__6183),
            .in2(N__6045),
            .in3(N__6630),
            .lcout(\display1.prescaler8_21 ),
            .ltout(\display1.prescaler8_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_0_LC_3_13_5 .C_ON=1'b0;
    defparam \display1.prescaler_0_LC_3_13_5 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_0_LC_3_13_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \display1.prescaler_0_LC_3_13_5  (
            .in0(N__6271),
            .in1(N__6226),
            .in2(N__6042),
            .in3(N__6148),
            .lcout(\display1.prescalerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14270),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_6_LC_3_13_6 .C_ON=1'b0;
    defparam \display1.prescaler_6_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_6_LC_3_13_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display1.prescaler_6_LC_3_13_6  (
            .in0(N__6308),
            .in1(N__6272),
            .in2(N__6233),
            .in3(N__6411),
            .lcout(\display1.prescalerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14270),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_1_LC_3_13_7 .C_ON=1'b0;
    defparam \display1.prescaler_1_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_1_LC_3_13_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \display1.prescaler_1_LC_3_13_7  (
            .in0(N__6167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6149),
            .lcout(\display1.prescalerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14270),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_9_LC_3_14_0 .C_ON=1'b0;
    defparam \display1.prescaler_9_LC_3_14_0 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_9_LC_3_14_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display1.prescaler_9_LC_3_14_0  (
            .in0(N__6312),
            .in1(N__6224),
            .in2(N__6278),
            .in3(N__6339),
            .lcout(\display1.prescalerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14266),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNI0V011_16_LC_3_14_2 .C_ON=1'b0;
    defparam \display1.prescaler_RNI0V011_16_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNI0V011_16_LC_3_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display1.prescaler_RNI0V011_16_LC_3_14_2  (
            .in0(N__6525),
            .in1(N__6543),
            .in2(N__6504),
            .in3(N__6147),
            .lcout(\display1.prescaler8_17 ),
            .ltout(\display1.prescaler8_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_14_LC_3_14_3 .C_ON=1'b0;
    defparam \display1.prescaler_14_LC_3_14_3 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_14_LC_3_14_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \display1.prescaler_14_LC_3_14_3  (
            .in0(N__6222),
            .in1(N__6588),
            .in2(N__6315),
            .in3(N__6310),
            .lcout(\display1.prescalerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14266),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_15_LC_3_14_4 .C_ON=1'b0;
    defparam \display1.prescaler_15_LC_3_14_4 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_15_LC_3_14_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display1.prescaler_15_LC_3_14_4  (
            .in0(N__6311),
            .in1(N__6223),
            .in2(N__6277),
            .in3(N__6555),
            .lcout(\display1.prescalerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14266),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNIBG671_19_LC_3_15_0 .C_ON=1'b0;
    defparam \display1.prescaler_RNIBG671_19_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNIBG671_19_LC_3_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display1.prescaler_RNIBG671_19_LC_3_15_0  (
            .in0(N__6444),
            .in1(N__6462),
            .in2(N__6726),
            .in3(N__6480),
            .lcout(\display1.prescaler8_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNI9TOE_2_LC_5_12_6 .C_ON=1'b0;
    defparam \display1.prescaler_RNI9TOE_2_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNI9TOE_2_LC_5_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display1.prescaler_RNI9TOE_2_LC_5_12_6  (
            .in0(N__6065),
            .in1(N__6125),
            .in2(N__6399),
            .in3(N__6110),
            .lcout(\display1.prescaler8_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_2_cry_1_c_LC_5_13_0 .C_ON=1'b1;
    defparam \display1.prescaler_2_cry_1_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_2_cry_1_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \display1.prescaler_2_cry_1_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__6171),
            .in2(N__6153),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\display1.prescaler_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_2_LC_5_13_1 .C_ON=1'b1;
    defparam \display1.prescaler_2_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_2_LC_5_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_2_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__6126),
            .in2(_gnd_net_),
            .in3(N__6114),
            .lcout(\display1.prescalerZ0Z_2 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_1 ),
            .carryout(\display1.prescaler_2_cry_2 ),
            .clk(N__14264),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_3_LC_5_13_2 .C_ON=1'b1;
    defparam \display1.prescaler_3_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_3_LC_5_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_3_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__6111),
            .in2(_gnd_net_),
            .in3(N__6099),
            .lcout(\display1.prescalerZ0Z_3 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_2 ),
            .carryout(\display1.prescaler_2_cry_3 ),
            .clk(N__14264),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_4_LC_5_13_3 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_4_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_4_LC_5_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_4_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__6096),
            .in2(_gnd_net_),
            .in3(N__6069),
            .lcout(\display1.prescaler_2_4 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_3 ),
            .carryout(\display1.prescaler_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_5_LC_5_13_4 .C_ON=1'b1;
    defparam \display1.prescaler_5_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_5_LC_5_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_5_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__6066),
            .in2(_gnd_net_),
            .in3(N__6054),
            .lcout(\display1.prescalerZ0Z_5 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_4 ),
            .carryout(\display1.prescaler_2_cry_5 ),
            .clk(N__14264),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_6_LC_5_13_5 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_6_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_6_LC_5_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_6_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__6426),
            .in2(_gnd_net_),
            .in3(N__6402),
            .lcout(\display1.prescaler_2_6 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_5 ),
            .carryout(\display1.prescaler_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_7_LC_5_13_6 .C_ON=1'b1;
    defparam \display1.prescaler_7_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_7_LC_5_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_7_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__6398),
            .in2(_gnd_net_),
            .in3(N__6384),
            .lcout(\display1.prescalerZ0Z_7 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_6 ),
            .carryout(\display1.prescaler_2_cry_7 ),
            .clk(N__14264),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_8_LC_5_13_7 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_8_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_8_LC_5_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_8_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__6381),
            .in2(_gnd_net_),
            .in3(N__6357),
            .lcout(\display1.prescaler_2_8 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_7 ),
            .carryout(\display1.prescaler_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_9_LC_5_14_0 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_9_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_9_LC_5_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_9_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__6354),
            .in2(_gnd_net_),
            .in3(N__6330),
            .lcout(\display1.prescaler_2_9 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\display1.prescaler_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_10_LC_5_14_1 .C_ON=1'b1;
    defparam \display1.prescaler_10_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_10_LC_5_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_10_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__6642),
            .in2(_gnd_net_),
            .in3(N__6327),
            .lcout(\display1.prescalerZ0Z_10 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_9 ),
            .carryout(\display1.prescaler_2_cry_10 ),
            .clk(N__14261),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_11_LC_5_14_2 .C_ON=1'b1;
    defparam \display1.prescaler_11_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_11_LC_5_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_11_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__6669),
            .in2(_gnd_net_),
            .in3(N__6324),
            .lcout(\display1.prescalerZ0Z_11 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_10 ),
            .carryout(\display1.prescaler_2_cry_11 ),
            .clk(N__14261),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_12_LC_5_14_3 .C_ON=1'b1;
    defparam \display1.prescaler_12_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_12_LC_5_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_12_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__6681),
            .in2(_gnd_net_),
            .in3(N__6321),
            .lcout(\display1.prescalerZ0Z_12 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_11 ),
            .carryout(\display1.prescaler_2_cry_12 ),
            .clk(N__14261),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_13_LC_5_14_4 .C_ON=1'b1;
    defparam \display1.prescaler_13_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_13_LC_5_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_13_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__6656),
            .in2(_gnd_net_),
            .in3(N__6318),
            .lcout(\display1.prescalerZ0Z_13 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_12 ),
            .carryout(\display1.prescaler_2_cry_13 ),
            .clk(N__14261),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_14_LC_5_14_5 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_14_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_14_LC_5_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_14_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__6603),
            .in2(_gnd_net_),
            .in3(N__6579),
            .lcout(\display1.prescaler_2_14 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_13 ),
            .carryout(\display1.prescaler_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNO_0_15_LC_5_14_6 .C_ON=1'b1;
    defparam \display1.prescaler_RNO_0_15_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNO_0_15_LC_5_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_RNO_0_15_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__6575),
            .in2(_gnd_net_),
            .in3(N__6546),
            .lcout(\display1.prescaler_2_15 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_14 ),
            .carryout(\display1.prescaler_2_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_16_LC_5_14_7 .C_ON=1'b1;
    defparam \display1.prescaler_16_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_16_LC_5_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_16_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__6542),
            .in2(_gnd_net_),
            .in3(N__6528),
            .lcout(\display1.prescalerZ0Z_16 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_15 ),
            .carryout(\display1.prescaler_2_cry_16 ),
            .clk(N__14261),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_17_LC_5_15_0 .C_ON=1'b1;
    defparam \display1.prescaler_17_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_17_LC_5_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_17_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__6524),
            .in2(_gnd_net_),
            .in3(N__6507),
            .lcout(\display1.prescalerZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\display1.prescaler_2_cry_17 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_18_LC_5_15_1 .C_ON=1'b1;
    defparam \display1.prescaler_18_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_18_LC_5_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_18_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__6497),
            .in2(_gnd_net_),
            .in3(N__6483),
            .lcout(\display1.prescalerZ0Z_18 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_17 ),
            .carryout(\display1.prescaler_2_cry_18 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_19_LC_5_15_2 .C_ON=1'b1;
    defparam \display1.prescaler_19_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_19_LC_5_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_19_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__6479),
            .in2(_gnd_net_),
            .in3(N__6465),
            .lcout(\display1.prescalerZ0Z_19 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_18 ),
            .carryout(\display1.prescaler_2_cry_19 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_20_LC_5_15_3 .C_ON=1'b1;
    defparam \display1.prescaler_20_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_20_LC_5_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_20_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__6461),
            .in2(_gnd_net_),
            .in3(N__6447),
            .lcout(\display1.prescalerZ0Z_20 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_19 ),
            .carryout(\display1.prescaler_2_cry_20 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_21_LC_5_15_4 .C_ON=1'b1;
    defparam \display1.prescaler_21_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_21_LC_5_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_21_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__6443),
            .in2(_gnd_net_),
            .in3(N__6429),
            .lcout(\display1.prescalerZ0Z_21 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_20 ),
            .carryout(\display1.prescaler_2_cry_21 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_22_LC_5_15_5 .C_ON=1'b1;
    defparam \display1.prescaler_22_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_22_LC_5_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display1.prescaler_22_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__6722),
            .in2(_gnd_net_),
            .in3(N__6708),
            .lcout(\display1.prescalerZ0Z_22 ),
            .ltout(),
            .carryin(\display1.prescaler_2_cry_21 ),
            .carryout(\display1.prescaler_2_cry_22 ),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_23_LC_5_15_6 .C_ON=1'b0;
    defparam \display1.prescaler_23_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \display1.prescaler_23_LC_5_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \display1.prescaler_23_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__6695),
            .in2(_gnd_net_),
            .in3(N__6705),
            .lcout(\display1.prescalerZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14258),
            .ce(),
            .sr(_gnd_net_));
    defparam \display1.prescaler_RNI24371_10_LC_5_15_7 .C_ON=1'b0;
    defparam \display1.prescaler_RNI24371_10_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \display1.prescaler_RNI24371_10_LC_5_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display1.prescaler_RNI24371_10_LC_5_15_7  (
            .in0(N__6680),
            .in1(N__6668),
            .in2(N__6657),
            .in3(N__6641),
            .lcout(\display1.prescaler8_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_RNIKI1C_LC_6_13_1 .C_ON=1'b0;
    defparam \d1.sync_1_RNIKI1C_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \d1.sync_1_RNIKI1C_LC_6_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \d1.sync_1_RNIKI1C_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__6944),
            .in2(_gnd_net_),
            .in3(N__9065),
            .lcout(\d1.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_stored_e_0_3_LC_6_14_0.C_ON=1'b0;
    defparam mins_stored_e_0_3_LC_6_14_0.SEQ_MODE=4'b1000;
    defparam mins_stored_e_0_3_LC_6_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 mins_stored_e_0_3_LC_6_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13899),
            .lcout(mins_storedZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14252),
            .ce(N__10774),
            .sr(_gnd_net_));
    defparam \d1.count_1_LC_6_15_0 .C_ON=1'b0;
    defparam \d1.count_1_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \d1.count_1_LC_6_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \d1.count_1_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__6917),
            .in2(_gnd_net_),
            .in3(N__8309),
            .lcout(\d1.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14245),
            .ce(),
            .sr(N__7071));
    defparam \d1.count_RNI0AFK_0_16_LC_6_16_1 .C_ON=1'b0;
    defparam \d1.count_RNI0AFK_0_16_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI0AFK_0_16_LC_6_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI0AFK_0_16_LC_6_16_1  (
            .in0(N__6913),
            .in1(N__7090),
            .in2(N__6894),
            .in3(N__7112),
            .lcout(\d1.g0_1_a5_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI0AFK_16_LC_6_16_6 .C_ON=1'b0;
    defparam \d1.count_RNI0AFK_16_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI0AFK_16_LC_6_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI0AFK_16_LC_6_16_6  (
            .in0(N__7111),
            .in1(N__6889),
            .in2(N__7092),
            .in3(N__6912),
            .lcout(\d1.trans_up_1_11 ),
            .ltout(\d1.trans_up_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIRPKB1_LC_6_16_7 .C_ON=1'b0;
    defparam \d1.state_RNIRPKB1_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIRPKB1_LC_6_16_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \d1.state_RNIRPKB1_LC_6_16_7  (
            .in0(N__9048),
            .in1(N__12798),
            .in2(N__6606),
            .in3(N__11902),
            .lcout(\d1.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.stateZ0_LC_6_17_4 .C_ON=1'b0;
    defparam \d1.stateZ0_LC_6_17_4 .SEQ_MODE=4'b1000;
    defparam \d1.stateZ0_LC_6_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d1.stateZ0_LC_6_17_4  (
            .in0(_gnd_net_),
            .in1(N__9052),
            .in2(_gnd_net_),
            .in3(N__10221),
            .lcout(\d1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14231),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNIQ0UE1_22_LC_7_11_1 .C_ON=1'b0;
    defparam \a.count_RNIQ0UE1_22_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \a.count_RNIQ0UE1_22_LC_7_11_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \a.count_RNIQ0UE1_22_LC_7_11_1  (
            .in0(N__7005),
            .in1(N__7020),
            .in2(N__7041),
            .in3(N__7524),
            .lcout(),
            .ltout(\a.BUZZER3_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNI7VOF2_4_LC_7_11_2 .C_ON=1'b0;
    defparam \a.count_RNI7VOF2_4_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \a.count_RNI7VOF2_4_LC_7_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \a.count_RNI7VOF2_4_LC_7_11_2  (
            .in0(N__10689),
            .in1(N__7281),
            .in2(N__6753),
            .in3(N__8662),
            .lcout(\a.BUZZER3_20 ),
            .ltout(\a.BUZZER3_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.BUZZER_LC_7_11_3 .C_ON=1'b0;
    defparam \a.BUZZER_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \a.BUZZER_LC_7_11_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \a.BUZZER_LC_7_11_3  (
            .in0(N__6737),
            .in1(N__6840),
            .in2(N__6750),
            .in3(N__6783),
            .lcout(BUZZER_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14262),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNI39TE1_10_LC_7_11_5 .C_ON=1'b0;
    defparam \a.count_RNI39TE1_10_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \a.count_RNI39TE1_10_LC_7_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \a.count_RNI39TE1_10_LC_7_11_5  (
            .in0(N__7236),
            .in1(N__7251),
            .in2(N__7179),
            .in3(N__7266),
            .lcout(\a.BUZZER3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_11_LC_7_12_0 .C_ON=1'b0;
    defparam \a.count_11_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \a.count_11_LC_7_12_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_11_LC_7_12_0  (
            .in0(N__6775),
            .in1(N__6863),
            .in2(N__6843),
            .in3(N__7140),
            .lcout(\a.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_10_LC_7_12_1 .C_ON=1'b0;
    defparam \a.count_10_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \a.count_10_LC_7_12_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_10_LC_7_12_1  (
            .in0(N__6862),
            .in1(N__6774),
            .in2(N__6841),
            .in3(N__7164),
            .lcout(\a.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_14_LC_7_12_2 .C_ON=1'b0;
    defparam \a.count_14_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \a.count_14_LC_7_12_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_14_LC_7_12_2  (
            .in0(N__6778),
            .in1(N__6866),
            .in2(N__6845),
            .in3(N__7344),
            .lcout(\a.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNIE4K61_11_LC_7_12_3 .C_ON=1'b0;
    defparam \a.count_RNIE4K61_11_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \a.count_RNIE4K61_11_LC_7_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \a.count_RNIE4K61_11_LC_7_12_3  (
            .in0(N__7376),
            .in1(N__7397),
            .in2(N__7155),
            .in3(N__7355),
            .lcout(\a.BUZZER3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_13_LC_7_12_4 .C_ON=1'b0;
    defparam \a.count_13_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \a.count_13_LC_7_12_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_13_LC_7_12_4  (
            .in0(N__6777),
            .in1(N__6865),
            .in2(N__6844),
            .in3(N__7365),
            .lcout(\a.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_8_LC_7_12_6 .C_ON=1'b0;
    defparam \a.count_8_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \a.count_8_LC_7_12_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_8_LC_7_12_6  (
            .in0(N__6779),
            .in1(N__6867),
            .in2(N__6846),
            .in3(N__7203),
            .lcout(\a.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_12_LC_7_12_7 .C_ON=1'b0;
    defparam \a.count_12_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \a.count_12_LC_7_12_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \a.count_12_LC_7_12_7  (
            .in0(N__6864),
            .in1(N__6776),
            .in2(N__6842),
            .in3(N__7386),
            .lcout(\a.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14259),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNIS97C1_23_LC_7_13_1 .C_ON=1'b0;
    defparam \a.count_RNIS97C1_23_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \a.count_RNIS97C1_23_LC_7_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \a.count_RNIS97C1_23_LC_7_13_1  (
            .in0(N__7505),
            .in1(N__7194),
            .in2(N__7221),
            .in3(N__7490),
            .lcout(\a.BUZZER3_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_LC_7_13_2 .C_ON=1'b0;
    defparam \d1.sync_1_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \d1.sync_1_LC_7_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d1.sync_1_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13917),
            .lcout(\d1.syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14253),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNISJL61_25_LC_7_13_3 .C_ON=1'b0;
    defparam \a.count_RNISJL61_25_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \a.count_RNISJL61_25_LC_7_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \a.count_RNISJL61_25_LC_7_13_3  (
            .in0(N__7334),
            .in1(N__7304),
            .in2(N__7473),
            .in3(N__7319),
            .lcout(),
            .ltout(\a.BUZZER3_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNIUI705_11_LC_7_13_4 .C_ON=1'b0;
    defparam \a.count_RNIUI705_11_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \a.count_RNIUI705_11_LC_7_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \a.count_RNIUI705_11_LC_7_13_4  (
            .in0(N__6798),
            .in1(N__6792),
            .in2(N__6786),
            .in3(N__7404),
            .lcout(\a.BUZZER3_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_LC_7_14_0.C_ON=1'b0;
    defparam prescaler_1_LC_7_14_0.SEQ_MODE=4'b1000;
    defparam prescaler_1_LC_7_14_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 prescaler_1_LC_7_14_0 (
            .in0(N__7676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7652),
            .lcout(prescalerZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14246),
            .ce(N__8053),
            .sr(_gnd_net_));
    defparam prescaler_0_LC_7_14_1.C_ON=1'b0;
    defparam prescaler_0_LC_7_14_1.SEQ_MODE=4'b1000;
    defparam prescaler_0_LC_7_14_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 prescaler_0_LC_7_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7675),
            .lcout(prescalerZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14246),
            .ce(N__8053),
            .sr(_gnd_net_));
    defparam \d1.count_RNI2PCE_0_3_LC_7_15_0 .C_ON=1'b0;
    defparam \d1.count_RNI2PCE_0_3_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI2PCE_0_3_LC_7_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI2PCE_0_3_LC_7_15_0  (
            .in0(N__11025),
            .in1(N__11052),
            .in2(N__11001),
            .in3(N__10968),
            .lcout(\d1.g0_1_a5_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI5QJP_11_LC_7_15_2 .C_ON=1'b0;
    defparam \d1.count_RNI5QJP_11_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI5QJP_11_LC_7_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI5QJP_11_LC_7_15_2  (
            .in0(N__8611),
            .in1(N__8270),
            .in2(N__9066),
            .in3(N__8303),
            .lcout(\d1.g0_1_a5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_0_LC_7_15_3 .C_ON=1'b0;
    defparam \d1.count_0_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \d1.count_0_LC_7_15_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \d1.count_0_LC_7_15_3  (
            .in0(N__8304),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\d1.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14238),
            .ce(),
            .sr(N__7072));
    defparam \d1.count_RNI2PCE_3_LC_7_15_4 .C_ON=1'b0;
    defparam \d1.count_RNI2PCE_3_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI2PCE_3_LC_7_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI2PCE_3_LC_7_15_4  (
            .in0(N__11026),
            .in1(N__11053),
            .in2(N__11002),
            .in3(N__10969),
            .lcout(\d1.trans_up_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_1_RNI5IAP_LC_7_15_5 .C_ON=1'b0;
    defparam \d1.sync_1_RNI5IAP_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \d1.sync_1_RNI5IAP_LC_7_15_5 .LUT_INIT=16'b0010100000000000;
    LogicCell40 \d1.sync_1_RNI5IAP_LC_7_15_5  (
            .in0(N__7131),
            .in1(N__9056),
            .in2(N__6948),
            .in3(N__6966),
            .lcout(\d1.trans_up_1_12 ),
            .ltout(\d1.trans_up_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI9D0D1_3_LC_7_15_6 .C_ON=1'b0;
    defparam \d1.count_RNI9D0D1_3_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI9D0D1_3_LC_7_15_6 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \d1.count_RNI9D0D1_3_LC_7_15_6  (
            .in0(N__9167),
            .in1(_gnd_net_),
            .in2(N__6930),
            .in3(N__8331),
            .lcout(),
            .ltout(\d1.g1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIINS67_LC_7_15_7 .C_ON=1'b0;
    defparam \d1.state_RNIINS67_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIINS67_LC_7_15_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \d1.state_RNIINS67_LC_7_15_7  (
            .in0(N__6927),
            .in1(N__10167),
            .in2(N__6921),
            .in3(N__9126),
            .lcout(\d1.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.un3_count_cry_1_c_LC_7_16_0 .C_ON=1'b1;
    defparam \d1.un3_count_cry_1_c_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \d1.un3_count_cry_1_c_LC_7_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d1.un3_count_cry_1_c_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__8308),
            .in2(N__6918),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\d1.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_2_LC_7_16_1 .C_ON=1'b1;
    defparam \d1.count_2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \d1.count_2_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_2_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__6893),
            .in2(_gnd_net_),
            .in3(N__6876),
            .lcout(\d1.countZ0Z_2 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_1 ),
            .carryout(\d1.un3_count_cry_2 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_3_LC_7_16_2 .C_ON=1'b1;
    defparam \d1.count_3_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \d1.count_3_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_3_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__10973),
            .in2(_gnd_net_),
            .in3(N__6873),
            .lcout(\d1.countZ0Z_3 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_2 ),
            .carryout(\d1.un3_count_cry_3 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_4_LC_7_16_3 .C_ON=1'b1;
    defparam \d1.count_4_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \d1.count_4_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_4_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__11030),
            .in2(_gnd_net_),
            .in3(N__6870),
            .lcout(\d1.countZ0Z_4 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_3 ),
            .carryout(\d1.un3_count_cry_4 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_5_LC_7_16_4 .C_ON=1'b1;
    defparam \d1.count_5_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \d1.count_5_LC_7_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_5_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__11057),
            .in2(_gnd_net_),
            .in3(N__6990),
            .lcout(\d1.countZ0Z_5 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_4 ),
            .carryout(\d1.un3_count_cry_5 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_6_LC_7_16_5 .C_ON=1'b1;
    defparam \d1.count_6_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \d1.count_6_LC_7_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_6_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__11006),
            .in2(_gnd_net_),
            .in3(N__6987),
            .lcout(\d1.countZ0Z_6 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_5 ),
            .carryout(\d1.un3_count_cry_6 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_7_LC_7_16_6 .C_ON=1'b1;
    defparam \d1.count_7_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \d1.count_7_LC_7_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_7_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__8876),
            .in2(_gnd_net_),
            .in3(N__6984),
            .lcout(\d1.countZ0Z_7 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_6 ),
            .carryout(\d1.un3_count_cry_7 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_8_LC_7_16_7 .C_ON=1'b1;
    defparam \d1.count_8_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \d1.count_8_LC_7_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_8_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__8929),
            .in2(_gnd_net_),
            .in3(N__6981),
            .lcout(\d1.countZ0Z_8 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_7 ),
            .carryout(\d1.un3_count_cry_8 ),
            .clk(N__14232),
            .ce(),
            .sr(N__7073));
    defparam \d1.count_9_LC_7_17_0 .C_ON=1'b1;
    defparam \d1.count_9_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \d1.count_9_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_9_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__8956),
            .in2(_gnd_net_),
            .in3(N__6978),
            .lcout(\d1.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\d1.un3_count_cry_9 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_10_LC_7_17_1 .C_ON=1'b1;
    defparam \d1.count_10_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \d1.count_10_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_10_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__8899),
            .in2(_gnd_net_),
            .in3(N__6975),
            .lcout(\d1.countZ0Z_10 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_9 ),
            .carryout(\d1.un3_count_cry_10 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_11_LC_7_17_2 .C_ON=1'b1;
    defparam \d1.count_11_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \d1.count_11_LC_7_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_11_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__8269),
            .in2(_gnd_net_),
            .in3(N__6972),
            .lcout(\d1.countZ0Z_11 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_10 ),
            .carryout(\d1.un3_count_cry_11 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_12_LC_7_17_3 .C_ON=1'b1;
    defparam \d1.count_12_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \d1.count_12_LC_7_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_12_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__8610),
            .in2(_gnd_net_),
            .in3(N__6969),
            .lcout(\d1.countZ0Z_12 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_11 ),
            .carryout(\d1.un3_count_cry_12 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_13_LC_7_17_4 .C_ON=1'b1;
    defparam \d1.count_13_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \d1.count_13_LC_7_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_13_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__6965),
            .in2(_gnd_net_),
            .in3(N__6951),
            .lcout(\d1.countZ0Z_13 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_12 ),
            .carryout(\d1.un3_count_cry_13 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_14_LC_7_17_5 .C_ON=1'b1;
    defparam \d1.count_14_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \d1.count_14_LC_7_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_14_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__7130),
            .in2(_gnd_net_),
            .in3(N__7116),
            .lcout(\d1.countZ0Z_14 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_13 ),
            .carryout(\d1.un3_count_cry_14 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_15_LC_7_17_6 .C_ON=1'b1;
    defparam \d1.count_15_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \d1.count_15_LC_7_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d1.count_15_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__7113),
            .in2(_gnd_net_),
            .in3(N__7098),
            .lcout(\d1.countZ0Z_15 ),
            .ltout(),
            .carryin(\d1.un3_count_cry_14 ),
            .carryout(\d1.un3_count_cry_15 ),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d1.count_16_LC_7_17_7 .C_ON=1'b0;
    defparam \d1.count_16_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \d1.count_16_LC_7_17_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d1.count_16_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__7091),
            .in2(_gnd_net_),
            .in3(N__7095),
            .lcout(\d1.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14224),
            .ce(),
            .sr(N__7074));
    defparam \d2.sync_0_LC_7_20_5 .C_ON=1'b0;
    defparam \d2.sync_0_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \d2.sync_0_LC_7_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \d2.sync_0_LC_7_20_5  (
            .in0(N__7056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\d2.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14210),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_1_LC_8_10_7 .C_ON=1'b0;
    defparam \a.count_1_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \a.count_1_LC_8_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \a.count_1_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__8664),
            .in2(_gnd_net_),
            .in3(N__7040),
            .lcout(\a.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14263),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_1_cry_1_c_LC_8_11_0 .C_ON=1'b1;
    defparam \a.count_1_cry_1_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \a.count_1_cry_1_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \a.count_1_cry_1_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__7036),
            .in2(N__8663),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\a.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_2_LC_8_11_1 .C_ON=1'b1;
    defparam \a.count_2_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \a.count_2_LC_8_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_2_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__7019),
            .in2(_gnd_net_),
            .in3(N__7008),
            .lcout(\a.countZ0Z_2 ),
            .ltout(),
            .carryin(\a.count_1_cry_1 ),
            .carryout(\a.count_1_cry_2 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_3_LC_8_11_2 .C_ON=1'b1;
    defparam \a.count_3_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \a.count_3_LC_8_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_3_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__7004),
            .in2(_gnd_net_),
            .in3(N__6993),
            .lcout(\a.countZ0Z_3 ),
            .ltout(),
            .carryin(\a.count_1_cry_2 ),
            .carryout(\a.count_1_cry_3 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_4_LC_8_11_3 .C_ON=1'b1;
    defparam \a.count_4_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \a.count_4_LC_8_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_4_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__7280),
            .in2(_gnd_net_),
            .in3(N__7269),
            .lcout(\a.countZ0Z_4 ),
            .ltout(),
            .carryin(\a.count_1_cry_3 ),
            .carryout(\a.count_1_cry_4 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_5_LC_8_11_4 .C_ON=1'b1;
    defparam \a.count_5_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \a.count_5_LC_8_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_5_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__7265),
            .in2(_gnd_net_),
            .in3(N__7254),
            .lcout(\a.countZ0Z_5 ),
            .ltout(),
            .carryin(\a.count_1_cry_4 ),
            .carryout(\a.count_1_cry_5 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_6_LC_8_11_5 .C_ON=1'b1;
    defparam \a.count_6_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \a.count_6_LC_8_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_6_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__7250),
            .in2(_gnd_net_),
            .in3(N__7239),
            .lcout(\a.countZ0Z_6 ),
            .ltout(),
            .carryin(\a.count_1_cry_5 ),
            .carryout(\a.count_1_cry_6 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_7_LC_8_11_6 .C_ON=1'b1;
    defparam \a.count_7_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \a.count_7_LC_8_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_7_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__7235),
            .in2(_gnd_net_),
            .in3(N__7224),
            .lcout(\a.countZ0Z_7 ),
            .ltout(),
            .carryin(\a.count_1_cry_6 ),
            .carryout(\a.count_1_cry_7 ),
            .clk(N__14260),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_8_LC_8_11_7 .C_ON=1'b1;
    defparam \a.count_RNO_0_8_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_8_LC_8_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_8_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__7214),
            .in2(_gnd_net_),
            .in3(N__7197),
            .lcout(\a.count_1_8 ),
            .ltout(),
            .carryin(\a.count_1_cry_7 ),
            .carryout(\a.count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_9_LC_8_12_0 .C_ON=1'b1;
    defparam \a.count_9_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \a.count_9_LC_8_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_9_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__7193),
            .in2(_gnd_net_),
            .in3(N__7182),
            .lcout(\a.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\a.count_1_cry_9 ),
            .clk(N__14254),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_10_LC_8_12_1 .C_ON=1'b1;
    defparam \a.count_RNO_0_10_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_10_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_10_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__7175),
            .in2(_gnd_net_),
            .in3(N__7158),
            .lcout(\a.count_1_10 ),
            .ltout(),
            .carryin(\a.count_1_cry_9 ),
            .carryout(\a.count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_11_LC_8_12_2 .C_ON=1'b1;
    defparam \a.count_RNO_0_11_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_11_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_11_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__7151),
            .in2(_gnd_net_),
            .in3(N__7134),
            .lcout(\a.count_1_11 ),
            .ltout(),
            .carryin(\a.count_1_cry_10 ),
            .carryout(\a.count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_12_LC_8_12_3 .C_ON=1'b1;
    defparam \a.count_RNO_0_12_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_12_LC_8_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_12_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__7398),
            .in2(_gnd_net_),
            .in3(N__7380),
            .lcout(\a.count_1_12 ),
            .ltout(),
            .carryin(\a.count_1_cry_11 ),
            .carryout(\a.count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_13_LC_8_12_4 .C_ON=1'b1;
    defparam \a.count_RNO_0_13_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_13_LC_8_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_13_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__7377),
            .in2(_gnd_net_),
            .in3(N__7359),
            .lcout(\a.count_1_13 ),
            .ltout(),
            .carryin(\a.count_1_cry_12 ),
            .carryout(\a.count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNO_0_14_LC_8_12_5 .C_ON=1'b1;
    defparam \a.count_RNO_0_14_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \a.count_RNO_0_14_LC_8_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_RNO_0_14_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__7356),
            .in2(_gnd_net_),
            .in3(N__7338),
            .lcout(\a.count_1_14 ),
            .ltout(),
            .carryin(\a.count_1_cry_13 ),
            .carryout(\a.count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_15_LC_8_12_6 .C_ON=1'b1;
    defparam \a.count_15_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \a.count_15_LC_8_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_15_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__7335),
            .in2(_gnd_net_),
            .in3(N__7323),
            .lcout(\a.countZ0Z_15 ),
            .ltout(),
            .carryin(\a.count_1_cry_14 ),
            .carryout(\a.count_1_cry_15 ),
            .clk(N__14254),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_16_LC_8_12_7 .C_ON=1'b1;
    defparam \a.count_16_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \a.count_16_LC_8_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_16_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__7320),
            .in2(_gnd_net_),
            .in3(N__7308),
            .lcout(\a.countZ0Z_16 ),
            .ltout(),
            .carryin(\a.count_1_cry_15 ),
            .carryout(\a.count_1_cry_16 ),
            .clk(N__14254),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_17_LC_8_13_0 .C_ON=1'b1;
    defparam \a.count_17_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \a.count_17_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_17_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__7305),
            .in2(_gnd_net_),
            .in3(N__7293),
            .lcout(\a.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\a.count_1_cry_17 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_18_LC_8_13_1 .C_ON=1'b1;
    defparam \a.count_18_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \a.count_18_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_18_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__7458),
            .in2(_gnd_net_),
            .in3(N__7290),
            .lcout(\a.countZ0Z_18 ),
            .ltout(),
            .carryin(\a.count_1_cry_17 ),
            .carryout(\a.count_1_cry_18 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_19_LC_8_13_2 .C_ON=1'b1;
    defparam \a.count_19_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \a.count_19_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_19_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__7416),
            .in2(_gnd_net_),
            .in3(N__7287),
            .lcout(\a.countZ0Z_19 ),
            .ltout(),
            .carryin(\a.count_1_cry_18 ),
            .carryout(\a.count_1_cry_19 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_20_LC_8_13_3 .C_ON=1'b1;
    defparam \a.count_20_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \a.count_20_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_20_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__7430),
            .in2(_gnd_net_),
            .in3(N__7284),
            .lcout(\a.countZ0Z_20 ),
            .ltout(),
            .carryin(\a.count_1_cry_19 ),
            .carryout(\a.count_1_cry_20 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_21_LC_8_13_4 .C_ON=1'b1;
    defparam \a.count_21_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \a.count_21_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_21_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__7445),
            .in2(_gnd_net_),
            .in3(N__7527),
            .lcout(\a.countZ0Z_21 ),
            .ltout(),
            .carryin(\a.count_1_cry_20 ),
            .carryout(\a.count_1_cry_21 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_22_LC_8_13_5 .C_ON=1'b1;
    defparam \a.count_22_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \a.count_22_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_22_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__7523),
            .in2(_gnd_net_),
            .in3(N__7509),
            .lcout(\a.countZ0Z_22 ),
            .ltout(),
            .carryin(\a.count_1_cry_21 ),
            .carryout(\a.count_1_cry_22 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_23_LC_8_13_6 .C_ON=1'b1;
    defparam \a.count_23_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \a.count_23_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_23_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__7506),
            .in2(_gnd_net_),
            .in3(N__7494),
            .lcout(\a.countZ0Z_23 ),
            .ltout(),
            .carryin(\a.count_1_cry_22 ),
            .carryout(\a.count_1_cry_23 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_24_LC_8_13_7 .C_ON=1'b1;
    defparam \a.count_24_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \a.count_24_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \a.count_24_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__7491),
            .in2(_gnd_net_),
            .in3(N__7479),
            .lcout(\a.countZ0Z_24 ),
            .ltout(),
            .carryin(\a.count_1_cry_23 ),
            .carryout(\a.count_1_cry_24 ),
            .clk(N__14247),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_25_LC_8_14_0 .C_ON=1'b0;
    defparam \a.count_25_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \a.count_25_LC_8_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \a.count_25_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__7472),
            .in2(_gnd_net_),
            .in3(N__7476),
            .lcout(\a.countZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14239),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_1_c_RNO_LC_8_14_1.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_1_c_RNO_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_1_c_RNO_LC_8_14_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 decrement_time_0_prescaler10_1_c_RNO_LC_8_14_1 (
            .in0(N__7562),
            .in1(N__7547),
            .in2(N__7581),
            .in3(N__7595),
            .lcout(decrement_time_0_prescaler10_1_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_0_c_RNO_LC_8_14_2.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_0_c_RNO_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_0_c_RNO_LC_8_14_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 decrement_time_0_prescaler10_0_c_RNO_LC_8_14_2 (
            .in0(N__7614),
            .in1(N__7632),
            .in2(N__7677),
            .in3(N__7648),
            .lcout(decrement_time_0_prescaler10_0_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_RNIOGM61_18_LC_8_14_7 .C_ON=1'b0;
    defparam \a.count_RNIOGM61_18_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \a.count_RNIOGM61_18_LC_8_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \a.count_RNIOGM61_18_LC_8_14_7  (
            .in0(N__7457),
            .in1(N__7446),
            .in2(N__7431),
            .in3(N__7415),
            .lcout(\a.BUZZER3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_1_c_LC_8_15_0.C_ON=1'b1;
    defparam prescaler_1_cry_1_c_LC_8_15_0.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_1_c_LC_8_15_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 prescaler_1_cry_1_c_LC_8_15_0 (
            .in0(_gnd_net_),
            .in1(N__7674),
            .in2(N__7653),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(prescaler_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_2_LC_8_15_1.C_ON=1'b1;
    defparam prescaler_2_LC_8_15_1.SEQ_MODE=4'b1000;
    defparam prescaler_2_LC_8_15_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_2_LC_8_15_1 (
            .in0(_gnd_net_),
            .in1(N__7631),
            .in2(_gnd_net_),
            .in3(N__7617),
            .lcout(prescalerZ0Z_2),
            .ltout(),
            .carryin(prescaler_1_cry_1),
            .carryout(prescaler_1_cry_2),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_3_LC_8_15_2.C_ON=1'b1;
    defparam prescaler_3_LC_8_15_2.SEQ_MODE=4'b1000;
    defparam prescaler_3_LC_8_15_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_3_LC_8_15_2 (
            .in0(_gnd_net_),
            .in1(N__7613),
            .in2(_gnd_net_),
            .in3(N__7599),
            .lcout(prescalerZ0Z_3),
            .ltout(),
            .carryin(prescaler_1_cry_2),
            .carryout(prescaler_1_cry_3),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_4_LC_8_15_3.C_ON=1'b1;
    defparam prescaler_4_LC_8_15_3.SEQ_MODE=4'b1000;
    defparam prescaler_4_LC_8_15_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_4_LC_8_15_3 (
            .in0(_gnd_net_),
            .in1(N__7596),
            .in2(_gnd_net_),
            .in3(N__7584),
            .lcout(prescalerZ0Z_4),
            .ltout(),
            .carryin(prescaler_1_cry_3),
            .carryout(prescaler_1_cry_4),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_5_LC_8_15_4.C_ON=1'b1;
    defparam prescaler_5_LC_8_15_4.SEQ_MODE=4'b1000;
    defparam prescaler_5_LC_8_15_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_5_LC_8_15_4 (
            .in0(_gnd_net_),
            .in1(N__7580),
            .in2(_gnd_net_),
            .in3(N__7566),
            .lcout(prescalerZ0Z_5),
            .ltout(),
            .carryin(prescaler_1_cry_4),
            .carryout(prescaler_1_cry_5),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_6_LC_8_15_5.C_ON=1'b1;
    defparam prescaler_6_LC_8_15_5.SEQ_MODE=4'b1000;
    defparam prescaler_6_LC_8_15_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_6_LC_8_15_5 (
            .in0(_gnd_net_),
            .in1(N__7563),
            .in2(_gnd_net_),
            .in3(N__7551),
            .lcout(prescalerZ0Z_6),
            .ltout(),
            .carryin(prescaler_1_cry_5),
            .carryout(prescaler_1_cry_6),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_7_LC_8_15_6.C_ON=1'b1;
    defparam prescaler_7_LC_8_15_6.SEQ_MODE=4'b1000;
    defparam prescaler_7_LC_8_15_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_7_LC_8_15_6 (
            .in0(_gnd_net_),
            .in1(N__7548),
            .in2(_gnd_net_),
            .in3(N__7536),
            .lcout(prescalerZ0Z_7),
            .ltout(),
            .carryin(prescaler_1_cry_6),
            .carryout(prescaler_1_cry_7),
            .clk(N__14233),
            .ce(N__8055),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_7_THRU_LUT4_0_LC_8_15_7.C_ON=1'b1;
    defparam prescaler_1_cry_7_THRU_LUT4_0_LC_8_15_7.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_7_THRU_LUT4_0_LC_8_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_7_THRU_LUT4_0_LC_8_15_7 (
            .in0(_gnd_net_),
            .in1(N__7902),
            .in2(_gnd_net_),
            .in3(N__7533),
            .lcout(prescaler_1_cry_7_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_7),
            .carryout(prescaler_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_9_LC_8_16_0.C_ON=1'b1;
    defparam prescaler_9_LC_8_16_0.SEQ_MODE=4'b1000;
    defparam prescaler_9_LC_8_16_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_9_LC_8_16_0 (
            .in0(_gnd_net_),
            .in1(N__8468),
            .in2(_gnd_net_),
            .in3(N__7530),
            .lcout(prescalerZ0Z_9),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(prescaler_1_cry_9),
            .clk(N__14225),
            .ce(N__8056),
            .sr(_gnd_net_));
    defparam prescaler_10_LC_8_16_1.C_ON=1'b1;
    defparam prescaler_10_LC_8_16_1.SEQ_MODE=4'b1000;
    defparam prescaler_10_LC_8_16_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_10_LC_8_16_1 (
            .in0(_gnd_net_),
            .in1(N__8495),
            .in2(_gnd_net_),
            .in3(N__7704),
            .lcout(prescalerZ0Z_10),
            .ltout(),
            .carryin(prescaler_1_cry_9),
            .carryout(prescaler_1_cry_10),
            .clk(N__14225),
            .ce(N__8056),
            .sr(_gnd_net_));
    defparam prescaler_11_LC_8_16_2.C_ON=1'b1;
    defparam prescaler_11_LC_8_16_2.SEQ_MODE=4'b1000;
    defparam prescaler_11_LC_8_16_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_11_LC_8_16_2 (
            .in0(_gnd_net_),
            .in1(N__8481),
            .in2(_gnd_net_),
            .in3(N__7701),
            .lcout(prescalerZ0Z_11),
            .ltout(),
            .carryin(prescaler_1_cry_10),
            .carryout(prescaler_1_cry_11),
            .clk(N__14225),
            .ce(N__8056),
            .sr(_gnd_net_));
    defparam prescaler_12_LC_8_16_3.C_ON=1'b1;
    defparam prescaler_12_LC_8_16_3.SEQ_MODE=4'b1000;
    defparam prescaler_12_LC_8_16_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_12_LC_8_16_3 (
            .in0(_gnd_net_),
            .in1(N__8454),
            .in2(_gnd_net_),
            .in3(N__7698),
            .lcout(prescalerZ0Z_12),
            .ltout(),
            .carryin(prescaler_1_cry_11),
            .carryout(prescaler_1_cry_12),
            .clk(N__14225),
            .ce(N__8056),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_12_THRU_LUT4_0_LC_8_16_4.C_ON=1'b1;
    defparam prescaler_1_cry_12_THRU_LUT4_0_LC_8_16_4.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_12_THRU_LUT4_0_LC_8_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_12_THRU_LUT4_0_LC_8_16_4 (
            .in0(_gnd_net_),
            .in1(N__8202),
            .in2(_gnd_net_),
            .in3(N__7695),
            .lcout(prescaler_1_cry_12_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_12),
            .carryout(prescaler_1_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_13_THRU_LUT4_0_LC_8_16_5.C_ON=1'b1;
    defparam prescaler_1_cry_13_THRU_LUT4_0_LC_8_16_5.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_13_THRU_LUT4_0_LC_8_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_13_THRU_LUT4_0_LC_8_16_5 (
            .in0(_gnd_net_),
            .in1(N__8163),
            .in2(_gnd_net_),
            .in3(N__7692),
            .lcout(prescaler_1_cry_13_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_13),
            .carryout(prescaler_1_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_14_THRU_LUT4_0_LC_8_16_6.C_ON=1'b1;
    defparam prescaler_1_cry_14_THRU_LUT4_0_LC_8_16_6.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_14_THRU_LUT4_0_LC_8_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_14_THRU_LUT4_0_LC_8_16_6 (
            .in0(_gnd_net_),
            .in1(N__8127),
            .in2(_gnd_net_),
            .in3(N__7689),
            .lcout(prescaler_1_cry_14_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_14),
            .carryout(prescaler_1_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_15_THRU_LUT4_0_LC_8_16_7.C_ON=1'b1;
    defparam prescaler_1_cry_15_THRU_LUT4_0_LC_8_16_7.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_15_THRU_LUT4_0_LC_8_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_15_THRU_LUT4_0_LC_8_16_7 (
            .in0(_gnd_net_),
            .in1(N__8094),
            .in2(_gnd_net_),
            .in3(N__7686),
            .lcout(prescaler_1_cry_15_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_15),
            .carryout(prescaler_1_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_17_LC_8_17_0.C_ON=1'b1;
    defparam prescaler_17_LC_8_17_0.SEQ_MODE=4'b1000;
    defparam prescaler_17_LC_8_17_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_17_LC_8_17_0 (
            .in0(_gnd_net_),
            .in1(N__8399),
            .in2(_gnd_net_),
            .in3(N__7683),
            .lcout(prescalerZ0Z_17),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(prescaler_1_cry_17),
            .clk(N__14219),
            .ce(N__8057),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_17_THRU_LUT4_0_LC_8_17_1.C_ON=1'b1;
    defparam prescaler_1_cry_17_THRU_LUT4_0_LC_8_17_1.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_17_THRU_LUT4_0_LC_8_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_17_THRU_LUT4_0_LC_8_17_1 (
            .in0(_gnd_net_),
            .in1(N__7953),
            .in2(_gnd_net_),
            .in3(N__7680),
            .lcout(prescaler_1_cry_17_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_17),
            .carryout(prescaler_1_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_19_LC_8_17_2.C_ON=1'b1;
    defparam prescaler_19_LC_8_17_2.SEQ_MODE=4'b1000;
    defparam prescaler_19_LC_8_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_19_LC_8_17_2 (
            .in0(_gnd_net_),
            .in1(N__8385),
            .in2(_gnd_net_),
            .in3(N__7731),
            .lcout(prescalerZ0Z_19),
            .ltout(),
            .carryin(prescaler_1_cry_18),
            .carryout(prescaler_1_cry_19),
            .clk(N__14219),
            .ce(N__8057),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_19_THRU_LUT4_0_LC_8_17_3.C_ON=1'b1;
    defparam prescaler_1_cry_19_THRU_LUT4_0_LC_8_17_3.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_19_THRU_LUT4_0_LC_8_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_19_THRU_LUT4_0_LC_8_17_3 (
            .in0(_gnd_net_),
            .in1(N__8031),
            .in2(_gnd_net_),
            .in3(N__7728),
            .lcout(prescaler_1_cry_19_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_19),
            .carryout(prescaler_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_20_THRU_LUT4_0_LC_8_17_4.C_ON=1'b1;
    defparam prescaler_1_cry_20_THRU_LUT4_0_LC_8_17_4.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_20_THRU_LUT4_0_LC_8_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_20_THRU_LUT4_0_LC_8_17_4 (
            .in0(_gnd_net_),
            .in1(N__8007),
            .in2(_gnd_net_),
            .in3(N__7725),
            .lcout(prescaler_1_cry_20_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_20),
            .carryout(prescaler_1_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_21_THRU_LUT4_0_LC_8_17_5.C_ON=1'b1;
    defparam prescaler_1_cry_21_THRU_LUT4_0_LC_8_17_5.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_21_THRU_LUT4_0_LC_8_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_21_THRU_LUT4_0_LC_8_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7983),
            .in3(N__7722),
            .lcout(prescaler_1_cry_21_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_21),
            .carryout(prescaler_1_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_22_THRU_LUT4_0_LC_8_17_6.C_ON=1'b1;
    defparam prescaler_1_cry_22_THRU_LUT4_0_LC_8_17_6.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_22_THRU_LUT4_0_LC_8_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_22_THRU_LUT4_0_LC_8_17_6 (
            .in0(_gnd_net_),
            .in1(N__7866),
            .in2(_gnd_net_),
            .in3(N__7719),
            .lcout(prescaler_1_cry_22_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_22),
            .carryout(prescaler_1_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_23_THRU_LUT4_0_LC_8_17_7.C_ON=1'b1;
    defparam prescaler_1_cry_23_THRU_LUT4_0_LC_8_17_7.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_23_THRU_LUT4_0_LC_8_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_23_THRU_LUT4_0_LC_8_17_7 (
            .in0(_gnd_net_),
            .in1(N__7833),
            .in2(_gnd_net_),
            .in3(N__7716),
            .lcout(prescaler_1_cry_23_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_23),
            .carryout(prescaler_1_cry_24),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_25_LC_8_18_0.C_ON=1'b1;
    defparam prescaler_25_LC_8_18_0.SEQ_MODE=4'b1000;
    defparam prescaler_25_LC_8_18_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescaler_25_LC_8_18_0 (
            .in0(_gnd_net_),
            .in1(N__8426),
            .in2(_gnd_net_),
            .in3(N__7713),
            .lcout(prescalerZ0Z_25),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(prescaler_1_cry_25),
            .clk(N__14215),
            .ce(N__8058),
            .sr(_gnd_net_));
    defparam prescaler_1_cry_25_THRU_LUT4_0_LC_8_18_1.C_ON=1'b1;
    defparam prescaler_1_cry_25_THRU_LUT4_0_LC_8_18_1.SEQ_MODE=4'b0000;
    defparam prescaler_1_cry_25_THRU_LUT4_0_LC_8_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescaler_1_cry_25_THRU_LUT4_0_LC_8_18_1 (
            .in0(_gnd_net_),
            .in1(N__7791),
            .in2(_gnd_net_),
            .in3(N__7710),
            .lcout(prescaler_1_cry_25_THRU_CO),
            .ltout(),
            .carryin(prescaler_1_cry_25),
            .carryout(prescaler_1_cry_26),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_27_LC_8_18_2.C_ON=1'b0;
    defparam prescaler_27_LC_8_18_2.SEQ_MODE=4'b1000;
    defparam prescaler_27_LC_8_18_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 prescaler_27_LC_8_18_2 (
            .in0(_gnd_net_),
            .in1(N__8412),
            .in2(_gnd_net_),
            .in3(N__7707),
            .lcout(prescalerZ0Z_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14215),
            .ce(N__8058),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_4_c_RNO_LC_9_11_0.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_4_c_RNO_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_4_c_RNO_LC_9_11_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 decrement_time_0_prescaler10_4_c_RNO_LC_9_11_0 (
            .in0(N__7891),
            .in1(N__7858),
            .in2(N__7829),
            .in3(N__7783),
            .lcout(decrement_time_0_prescaler10_4_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_8_LC_9_11_1.C_ON=1'b0;
    defparam prescaler_8_LC_9_11_1.SEQ_MODE=4'b1000;
    defparam prescaler_8_LC_9_11_1.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_8_LC_9_11_1 (
            .in0(N__7901),
            .in1(N__7914),
            .in2(_gnd_net_),
            .in3(N__9944),
            .lcout(prescalerZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_23_LC_9_11_2.C_ON=1'b0;
    defparam prescaler_23_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam prescaler_23_LC_9_11_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescaler_23_LC_9_11_2 (
            .in0(N__9941),
            .in1(N__7878),
            .in2(_gnd_net_),
            .in3(N__7859),
            .lcout(prescalerZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_24_LC_9_11_3.C_ON=1'b0;
    defparam prescaler_24_LC_9_11_3.SEQ_MODE=4'b1000;
    defparam prescaler_24_LC_9_11_3.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_24_LC_9_11_3 (
            .in0(N__7828),
            .in1(N__7845),
            .in2(_gnd_net_),
            .in3(N__9942),
            .lcout(prescalerZ0Z_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_26_LC_9_11_4.C_ON=1'b0;
    defparam prescaler_26_LC_9_11_4.SEQ_MODE=4'b1000;
    defparam prescaler_26_LC_9_11_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescaler_26_LC_9_11_4 (
            .in0(N__9943),
            .in1(N__7806),
            .in2(_gnd_net_),
            .in3(N__7784),
            .lcout(prescalerZ0Z_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_20_LC_9_11_5.C_ON=1'b0;
    defparam prescaler_20_LC_9_11_5.SEQ_MODE=4'b1000;
    defparam prescaler_20_LC_9_11_5.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_20_LC_9_11_5 (
            .in0(N__7770),
            .in1(N__8027),
            .in2(_gnd_net_),
            .in3(N__9938),
            .lcout(prescalerZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_21_LC_9_11_6.C_ON=1'b0;
    defparam prescaler_21_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam prescaler_21_LC_9_11_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescaler_21_LC_9_11_6 (
            .in0(N__9939),
            .in1(N__7755),
            .in2(_gnd_net_),
            .in3(N__8003),
            .lcout(prescalerZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam prescaler_22_LC_9_11_7.C_ON=1'b0;
    defparam prescaler_22_LC_9_11_7.SEQ_MODE=4'b1000;
    defparam prescaler_22_LC_9_11_7.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_22_LC_9_11_7 (
            .in0(N__7743),
            .in1(N__7972),
            .in2(_gnd_net_),
            .in3(N__9940),
            .lcout(prescalerZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14255),
            .ce(N__8052),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_2_c_RNO_LC_9_12_1.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_2_c_RNO_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_2_c_RNO_LC_9_12_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 decrement_time_0_prescaler10_2_c_RNO_LC_9_12_1 (
            .in0(N__8083),
            .in1(N__8119),
            .in2(N__8198),
            .in3(N__8155),
            .lcout(decrement_time_0_prescaler10_2_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescaler_13_LC_9_12_2.C_ON=1'b0;
    defparam prescaler_13_LC_9_12_2.SEQ_MODE=4'b1000;
    defparam prescaler_13_LC_9_12_2.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_13_LC_9_12_2 (
            .in0(N__8197),
            .in1(N__8214),
            .in2(_gnd_net_),
            .in3(N__9915),
            .lcout(prescalerZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14248),
            .ce(N__8054),
            .sr(_gnd_net_));
    defparam prescaler_14_LC_9_12_3.C_ON=1'b0;
    defparam prescaler_14_LC_9_12_3.SEQ_MODE=4'b1000;
    defparam prescaler_14_LC_9_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescaler_14_LC_9_12_3 (
            .in0(N__9916),
            .in1(N__8175),
            .in2(_gnd_net_),
            .in3(N__8156),
            .lcout(prescalerZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14248),
            .ce(N__8054),
            .sr(_gnd_net_));
    defparam prescaler_15_LC_9_12_4.C_ON=1'b0;
    defparam prescaler_15_LC_9_12_4.SEQ_MODE=4'b1000;
    defparam prescaler_15_LC_9_12_4.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_15_LC_9_12_4 (
            .in0(N__8120),
            .in1(N__8142),
            .in2(_gnd_net_),
            .in3(N__9917),
            .lcout(prescalerZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14248),
            .ce(N__8054),
            .sr(_gnd_net_));
    defparam prescaler_16_LC_9_12_5.C_ON=1'b0;
    defparam prescaler_16_LC_9_12_5.SEQ_MODE=4'b1000;
    defparam prescaler_16_LC_9_12_5.LUT_INIT=16'b0001010000010100;
    LogicCell40 prescaler_16_LC_9_12_5 (
            .in0(N__9918),
            .in1(N__8106),
            .in2(N__8090),
            .in3(_gnd_net_),
            .lcout(prescalerZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14248),
            .ce(N__8054),
            .sr(_gnd_net_));
    defparam prescaler_18_LC_9_12_6.C_ON=1'b0;
    defparam prescaler_18_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam prescaler_18_LC_9_12_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 prescaler_18_LC_9_12_6 (
            .in0(N__7946),
            .in1(N__8070),
            .in2(_gnd_net_),
            .in3(N__9919),
            .lcout(prescalerZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14248),
            .ce(N__8054),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_3_c_RNO_LC_9_12_7.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_3_c_RNO_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_3_c_RNO_LC_9_12_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 decrement_time_0_prescaler10_3_c_RNO_LC_9_12_7 (
            .in0(N__8023),
            .in1(N__7999),
            .in2(N__7979),
            .in3(N__7945),
            .lcout(decrement_time_0_prescaler10_3_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_0_c_LC_9_13_0.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_0_c_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_0_c_LC_9_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_0_c_LC_9_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(decrement_time_0_prescaler10_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_1_c_LC_9_13_1.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_1_c_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_1_c_LC_9_13_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_1_c_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7923),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_0),
            .carryout(decrement_time_0_prescaler10_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_2_c_LC_9_13_2.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_2_c_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_2_c_LC_9_13_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_2_c_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_1),
            .carryout(decrement_time_0_prescaler10_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_3_c_LC_9_13_3.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_3_c_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_3_c_LC_9_13_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_3_c_LC_9_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8238),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_2),
            .carryout(decrement_time_0_prescaler10_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_4_c_LC_9_13_4.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_4_c_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_4_c_LC_9_13_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_4_c_LC_9_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8229),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_3),
            .carryout(decrement_time_0_prescaler10_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_5_c_LC_9_13_5.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_5_c_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_5_c_LC_9_13_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_5_c_LC_9_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8442),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_4),
            .carryout(decrement_time_0_prescaler10_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_6_c_LC_9_13_6.C_ON=1'b1;
    defparam decrement_time_0_prescaler10_6_c_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_6_c_LC_9_13_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 decrement_time_0_prescaler10_6_c_LC_9_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8373),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(decrement_time_0_prescaler10_5),
            .carryout(decrement_time_0_prescaler10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_THRU_LUT4_0_LC_9_13_7.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_THRU_LUT4_0_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_THRU_LUT4_0_LC_9_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 decrement_time_0_prescaler10_THRU_LUT4_0_LC_9_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8217),
            .lcout(decrement_time_0_prescaler10_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_stored_e_0_0_LC_9_14_2.C_ON=1'b0;
    defparam mins_stored_e_0_0_LC_9_14_2.SEQ_MODE=4'b1000;
    defparam mins_stored_e_0_0_LC_9_14_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 mins_stored_e_0_0_LC_9_14_2 (
            .in0(N__13549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(mins_storedZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14234),
            .ce(N__10778),
            .sr(_gnd_net_));
    defparam mins_stored_e_0_1_LC_9_14_3.C_ON=1'b0;
    defparam mins_stored_e_0_1_LC_9_14_3.SEQ_MODE=4'b1000;
    defparam mins_stored_e_0_1_LC_9_14_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 mins_stored_e_0_1_LC_9_14_3 (
            .in0(N__13633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(mins_storedZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14234),
            .ce(N__10778),
            .sr(_gnd_net_));
    defparam mins_stored_e_0_2_LC_9_14_4.C_ON=1'b0;
    defparam mins_stored_e_0_2_LC_9_14_4.SEQ_MODE=4'b1000;
    defparam mins_stored_e_0_2_LC_9_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 mins_stored_e_0_2_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13788),
            .lcout(mins_storedZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14234),
            .ce(N__10778),
            .sr(_gnd_net_));
    defparam \d3.count_RNI1N275_12_LC_9_14_7 .C_ON=1'b0;
    defparam \d3.count_RNI1N275_12_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNI1N275_12_LC_9_14_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \d3.count_RNI1N275_12_LC_9_14_7  (
            .in0(N__8727),
            .in1(N__8706),
            .in2(N__9699),
            .in3(N__8628),
            .lcout(d3_trans_up_1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_6_LC_9_15_1 .C_ON=1'b0;
    defparam \d1.g0_6_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \d1.g0_6_LC_9_15_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \d1.g0_6_LC_9_15_1  (
            .in0(N__13544),
            .in1(N__13885),
            .in2(N__13646),
            .in3(N__13756),
            .lcout(),
            .ltout(\d1.mins27_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_0_LC_9_15_2 .C_ON=1'b0;
    defparam \d1.g2_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \d1.g2_0_LC_9_15_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \d1.g2_0_LC_9_15_2  (
            .in0(N__12114),
            .in1(N__11124),
            .in2(N__8355),
            .in3(N__8508),
            .lcout(),
            .ltout(\d1.g2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_0_o3_LC_9_15_3 .C_ON=1'b0;
    defparam \d1.g0_0_o3_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \d1.g0_0_o3_LC_9_15_3 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \d1.g0_0_o3_LC_9_15_3  (
            .in0(N__10494),
            .in1(N__8322),
            .in2(N__8352),
            .in3(N__10024),
            .lcout(\d1.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ten_secs_2_LC_9_15_4.C_ON=1'b0;
    defparam ten_secs_2_LC_9_15_4.SEQ_MODE=4'b1000;
    defparam ten_secs_2_LC_9_15_4.LUT_INIT=16'b0010100010001000;
    LogicCell40 ten_secs_2_LC_9_15_4 (
            .in0(N__10896),
            .in1(N__10589),
            .in2(N__12390),
            .in3(N__8747),
            .lcout(ten_secsZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14226),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI5FPI2_3_LC_9_15_5 .C_ON=1'b0;
    defparam \d1.count_RNI5FPI2_3_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI5FPI2_3_LC_9_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI5FPI2_3_LC_9_15_5  (
            .in0(N__8349),
            .in1(N__8340),
            .in2(N__10945),
            .in3(N__8850),
            .lcout(\d1.g0_1_a5_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_11_LC_9_15_6 .C_ON=1'b0;
    defparam \d1.g0_11_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \d1.g0_11_LC_9_15_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \d1.g0_11_LC_9_15_6  (
            .in0(N__13757),
            .in1(N__13614),
            .in2(N__13897),
            .in3(N__13545),
            .lcout(\d1.g0_0_0_a4_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_LC_9_15_7 .C_ON=1'b0;
    defparam \d1.g2_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_LC_9_15_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \d1.g2_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__11084),
            .in2(_gnd_net_),
            .in3(N__9816),
            .lcout(\d1.gZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIH1EH_7_LC_9_16_0 .C_ON=1'b0;
    defparam \d1.count_RNIH1EH_7_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIH1EH_7_LC_9_16_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.count_RNIH1EH_7_LC_9_16_0  (
            .in0(N__8933),
            .in1(N__8315),
            .in2(N__8280),
            .in3(N__8875),
            .lcout(\d1.g1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIQ6A21_11_LC_9_16_1 .C_ON=1'b0;
    defparam \d1.count_RNIQ6A21_11_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIQ6A21_11_LC_9_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNIQ6A21_11_LC_9_16_1  (
            .in0(N__8316),
            .in1(N__8276),
            .in2(N__8619),
            .in3(N__8849),
            .lcout(\d1.trans_up_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ten_secs_0_LC_9_16_2.C_ON=1'b0;
    defparam ten_secs_0_LC_9_16_2.SEQ_MODE=4'b1000;
    defparam ten_secs_0_LC_9_16_2.LUT_INIT=16'b0010001010001000;
    LogicCell40 ten_secs_0_LC_9_16_2 (
            .in0(N__10901),
            .in1(N__12429),
            .in2(_gnd_net_),
            .in3(N__8748),
            .lcout(ten_secsZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14220),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_2_LC_9_16_3 .C_ON=1'b0;
    defparam \d1.g2_2_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \d1.g2_2_LC_9_16_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \d1.g2_2_LC_9_16_3  (
            .in0(N__11710),
            .in1(N__11284),
            .in2(N__12799),
            .in3(N__9237),
            .lcout(\d1.g2_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.sync_1_LC_9_16_4 .C_ON=1'b0;
    defparam \d3.sync_1_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \d3.sync_1_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d3.sync_1_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8562),
            .lcout(\d3.syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14220),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_12_LC_9_16_6 .C_ON=1'b0;
    defparam \d1.g2_12_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \d1.g2_12_LC_9_16_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \d1.g2_12_LC_9_16_6  (
            .in0(N__12109),
            .in1(N__9258),
            .in2(N__12800),
            .in3(N__12356),
            .lcout(),
            .ltout(\d1.g2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_0_4_LC_9_16_7 .C_ON=1'b0;
    defparam \d1.g2_0_4_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_0_4_LC_9_16_7 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \d1.g2_0_4_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__8550),
            .in2(N__8502),
            .in3(N__11285),
            .lcout(\d1.g2_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_5_c_RNO_LC_9_17_0.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_5_c_RNO_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_5_c_RNO_LC_9_17_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 decrement_time_0_prescaler10_5_c_RNO_LC_9_17_0 (
            .in0(N__8499),
            .in1(N__8480),
            .in2(N__8469),
            .in3(N__8453),
            .lcout(decrement_time_0_prescaler10_5_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam decrement_time_0_prescaler10_6_c_RNO_LC_9_17_1.C_ON=1'b0;
    defparam decrement_time_0_prescaler10_6_c_RNO_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam decrement_time_0_prescaler10_6_c_RNO_LC_9_17_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 decrement_time_0_prescaler10_6_c_RNO_LC_9_17_1 (
            .in0(N__8427),
            .in1(N__8411),
            .in2(N__8400),
            .in3(N__8384),
            .lcout(decrement_time_0_prescaler10_6_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_15_LC_9_17_3 .C_ON=1'b0;
    defparam \d1.g2_15_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \d1.g2_15_LC_9_17_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_15_LC_9_17_3  (
            .in0(N__11493),
            .in1(N__11634),
            .in2(N__11712),
            .in3(N__11440),
            .lcout(),
            .ltout(\d1.g2_7_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_11_LC_9_17_4 .C_ON=1'b0;
    defparam \d1.g2_11_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \d1.g2_11_LC_9_17_4 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \d1.g2_11_LC_9_17_4  (
            .in0(N__11237),
            .in1(N__11180),
            .in2(N__8358),
            .in3(N__11903),
            .lcout(\d1.g2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNID2KP_9_LC_9_17_7 .C_ON=1'b0;
    defparam \d1.count_RNID2KP_9_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNID2KP_9_LC_9_17_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.count_RNID2KP_9_LC_9_17_7  (
            .in0(N__8612),
            .in1(N__8903),
            .in2(N__9076),
            .in3(N__8960),
            .lcout(\d1.g1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIVLG6B_LC_9_18_4 .C_ON=1'b0;
    defparam \d1.state_RNIVLG6B_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIVLG6B_LC_9_18_4 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \d1.state_RNIVLG6B_LC_9_18_4  (
            .in0(N__11541),
            .in1(N__10161),
            .in2(N__10188),
            .in3(N__10124),
            .lcout(\d1.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.sync_0_LC_9_18_5 .C_ON=1'b0;
    defparam \d3.sync_0_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \d3.sync_0_LC_9_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d3.sync_0_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8580),
            .lcout(\d3.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14211),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_5_LC_9_18_6 .C_ON=1'b0;
    defparam \d1.g2_5_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \d1.g2_5_LC_9_18_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_5_LC_9_18_6  (
            .in0(N__11492),
            .in1(N__11622),
            .in2(N__11711),
            .in3(N__11434),
            .lcout(\d1.g2_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_LC_9_18_7 .C_ON=1'b0;
    defparam \d2.sync_1_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \d2.sync_1_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d2.sync_1_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8541),
            .lcout(d2_sync_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14211),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_1_LC_9_19_3 .C_ON=1'b0;
    defparam \d2.count_1_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \d2.count_1_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \d2.count_1_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__11626),
            .in2(_gnd_net_),
            .in3(N__11439),
            .lcout(d2_count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14207),
            .ce(),
            .sr(N__10290));
    defparam \d2.count_0_LC_9_19_7 .C_ON=1'b0;
    defparam \d2.count_0_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_0_LC_9_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \d2.count_0_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11438),
            .lcout(d2_count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14207),
            .ce(),
            .sr(N__10290));
    defparam \d4.sync_1_LC_10_5_1 .C_ON=1'b0;
    defparam \d4.sync_1_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \d4.sync_1_LC_10_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d4.sync_1_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13311),
            .lcout(\d4.syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14271),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.sync_1_RNIQPEK_LC_10_8_7 .C_ON=1'b0;
    defparam \d4.sync_1_RNIQPEK_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \d4.sync_1_RNIQPEK_LC_10_8_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \d4.sync_1_RNIQPEK_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__8721),
            .in2(_gnd_net_),
            .in3(N__8795),
            .lcout(\d4.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_1_LC_10_10_0 .C_ON=1'b0;
    defparam \d4.count_1_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \d4.count_1_LC_10_10_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \d4.count_1_LC_10_10_0  (
            .in0(N__9362),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9337),
            .lcout(\d4.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14256),
            .ce(),
            .sr(N__9619));
    defparam \d4.count_0_LC_10_10_1 .C_ON=1'b0;
    defparam \d4.count_0_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \d4.count_0_LC_10_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \d4.count_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9361),
            .lcout(\d4.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14256),
            .ce(),
            .sr(N__9619));
    defparam \d1.g2_9_LC_10_11_0 .C_ON=1'b0;
    defparam \d1.g2_9_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \d1.g2_9_LC_10_11_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \d1.g2_9_LC_10_11_0  (
            .in0(N__13780),
            .in1(N__13671),
            .in2(N__13547),
            .in3(N__13898),
            .lcout(),
            .ltout(\d1.g2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_0_3_LC_10_11_1 .C_ON=1'b0;
    defparam \d1.g2_0_3_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \d1.g2_0_3_LC_10_11_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \d1.g2_0_3_LC_10_11_1  (
            .in0(N__11882),
            .in1(N__11238),
            .in2(N__8670),
            .in3(N__11181),
            .lcout(\d1.g2_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.ten_secs_1_sqmuxa_0_x1_LC_10_11_2 .C_ON=1'b0;
    defparam \d1.ten_secs_1_sqmuxa_0_x1_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \d1.ten_secs_1_sqmuxa_0_x1_LC_10_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \d1.ten_secs_1_sqmuxa_0_x1_LC_10_11_2  (
            .in0(N__12494),
            .in1(N__12449),
            .in2(N__10607),
            .in3(N__11881),
            .lcout(),
            .ltout(\d1.ten_secs_1_sqmuxa_0_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.ten_secs_1_sqmuxa_0_ns_LC_10_11_3 .C_ON=1'b0;
    defparam \d1.ten_secs_1_sqmuxa_0_ns_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \d1.ten_secs_1_sqmuxa_0_ns_LC_10_11_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \d1.ten_secs_1_sqmuxa_0_ns_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8667),
            .in3(N__12759),
            .lcout(\d1.ten_secs_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \a.count_0_LC_10_11_4 .C_ON=1'b0;
    defparam \a.count_0_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \a.count_0_LC_10_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \a.count_0_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8655),
            .lcout(\a.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14249),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_RNI5PSB_10_LC_10_11_5 .C_ON=1'b0;
    defparam \d4.count_RNI5PSB_10_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \d4.count_RNI5PSB_10_LC_10_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d4.count_RNI5PSB_10_LC_10_11_5  (
            .in0(N__9467),
            .in1(N__9452),
            .in2(N__9438),
            .in3(N__9482),
            .lcout(\d4.trans_up_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_RNIS9LE1_10_LC_10_12_1 .C_ON=1'b0;
    defparam \d3.count_RNIS9LE1_10_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNIS9LE1_10_LC_10_12_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d3.count_RNIS9LE1_10_LC_10_12_1  (
            .in0(N__9738),
            .in1(N__9580),
            .in2(N__9720),
            .in3(N__9603),
            .lcout(\d3.trans_up_1_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_1_LC_10_12_2 .C_ON=1'b0;
    defparam \d3.count_1_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \d3.count_1_LC_10_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \d3.count_1_LC_10_12_2  (
            .in0(N__9605),
            .in1(_gnd_net_),
            .in2(N__9587),
            .in3(_gnd_net_),
            .lcout(\d3.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14240),
            .ce(),
            .sr(N__9958));
    defparam \d3.count_0_LC_10_12_3 .C_ON=1'b0;
    defparam \d3.count_0_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \d3.count_0_LC_10_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \d3.count_0_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9604),
            .lcout(\d3.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14240),
            .ce(),
            .sr(N__9958));
    defparam \d4.count_RNICSOB_16_LC_10_12_4 .C_ON=1'b0;
    defparam \d4.count_RNICSOB_16_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \d4.count_RNICSOB_16_LC_10_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d4.count_RNICSOB_16_LC_10_12_4  (
            .in0(N__9653),
            .in1(N__9314),
            .in2(N__9636),
            .in3(N__9338),
            .lcout(\d4.trans_up_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_RNIE50C_3_LC_10_12_5 .C_ON=1'b0;
    defparam \d4.count_RNIE50C_3_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \d4.count_RNIE50C_3_LC_10_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d4.count_RNIE50C_3_LC_10_12_5  (
            .in0(N__9284),
            .in1(N__9269),
            .in2(N__9501),
            .in3(N__9299),
            .lcout(\d4.trans_up_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_RNIMDFN1_6_LC_10_13_0 .C_ON=1'b0;
    defparam \d3.count_RNIMDFN1_6_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNIMDFN1_6_LC_10_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d3.count_RNIMDFN1_6_LC_10_13_0  (
            .in0(N__9770),
            .in1(N__9785),
            .in2(N__9756),
            .in3(N__9800),
            .lcout(\d3.trans_up_1_15_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.sync_1_RNIHL7Q_LC_10_13_1 .C_ON=1'b0;
    defparam \d4.sync_1_RNIHL7Q_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \d4.sync_1_RNIHL7Q_LC_10_13_1 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \d4.sync_1_RNIHL7Q_LC_10_13_1  (
            .in0(N__9386),
            .in1(N__8720),
            .in2(N__9672),
            .in3(N__8792),
            .lcout(\d4.trans_up_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_RNI6TEN1_2_LC_10_13_2 .C_ON=1'b0;
    defparam \d3.count_RNI6TEN1_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNI6TEN1_2_LC_10_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d3.count_RNI6TEN1_2_LC_10_13_2  (
            .in0(N__9536),
            .in1(N__9551),
            .in2(N__9522),
            .in3(N__9566),
            .lcout(\d3.trans_up_1_15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.state_LC_10_13_3 .C_ON=1'b0;
    defparam \d4.state_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \d4.state_LC_10_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d4.state_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__8763),
            .in2(_gnd_net_),
            .in3(N__8794),
            .lcout(d4_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14235),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_RNIFDLK_11_LC_10_13_4 .C_ON=1'b0;
    defparam \d4.count_RNIFDLK_11_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \d4.count_RNIFDLK_11_LC_10_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d4.count_RNIFDLK_11_LC_10_13_4  (
            .in0(N__9419),
            .in1(N__9366),
            .in2(N__9405),
            .in3(N__8700),
            .lcout(),
            .ltout(\d4.trans_up_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_RNIQ4M62_11_LC_10_13_5 .C_ON=1'b0;
    defparam \d4.count_RNIQ4M62_11_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \d4.count_RNIQ4M62_11_LC_10_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d4.count_RNIQ4M62_11_LC_10_13_5  (
            .in0(N__8691),
            .in1(N__8685),
            .in2(N__8679),
            .in3(N__8676),
            .lcout(d4_trans_up_1),
            .ltout(d4_trans_up_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_1_sqmuxa_LC_10_13_6 .C_ON=1'b0;
    defparam \d1.state_1_sqmuxa_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \d1.state_1_sqmuxa_LC_10_13_6 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \d1.state_1_sqmuxa_LC_10_13_6  (
            .in0(N__8793),
            .in1(_gnd_net_),
            .in2(N__8808),
            .in3(N__9865),
            .lcout(\d1.state_1_sqmuxaZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ten_secs_RNO_0_1_LC_10_14_0.C_ON=1'b0;
    defparam ten_secs_RNO_0_1_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam ten_secs_RNO_0_1_LC_10_14_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 ten_secs_RNO_0_1_LC_10_14_0 (
            .in0(N__12436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8743),
            .lcout(),
            .ltout(ten_secs_r_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ten_secs_1_LC_10_14_1.C_ON=1'b0;
    defparam ten_secs_1_LC_10_14_1.SEQ_MODE=4'b1000;
    defparam ten_secs_1_LC_10_14_1.LUT_INIT=16'b0000000000101000;
    LogicCell40 ten_secs_1_LC_10_14_1 (
            .in0(N__10902),
            .in1(N__12490),
            .in2(N__8805),
            .in3(N__10825),
            .lcout(ten_secsZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14227),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_RNIEJS51_16_LC_10_14_2 .C_ON=1'b0;
    defparam \d3.count_RNIEJS51_16_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNIEJS51_16_LC_10_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d3.count_RNIEJS51_16_LC_10_14_2  (
            .in0(N__10666),
            .in1(N__10649),
            .in2(N__9837),
            .in3(N__10631),
            .lcout(\d3.trans_up_1_14_2 ),
            .ltout(\d3.trans_up_1_14_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.state_RNI7N9P6_LC_10_14_3 .C_ON=1'b0;
    defparam \d3.state_RNI7N9P6_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \d3.state_RNI7N9P6_LC_10_14_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \d3.state_RNI7N9P6_LC_10_14_3  (
            .in0(N__12576),
            .in1(N__12609),
            .in2(N__8802),
            .in3(N__11083),
            .lcout(s_cancel),
            .ltout(s_cancel_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.alarm_on_0_sqmuxa_LC_10_14_4 .C_ON=1'b0;
    defparam \d1.alarm_on_0_sqmuxa_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \d1.alarm_on_0_sqmuxa_LC_10_14_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \d1.alarm_on_0_sqmuxa_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__12770),
            .in2(N__8799),
            .in3(N__11886),
            .lcout(alarm_on_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.mins_stored_0_sqmuxa_LC_10_14_5 .C_ON=1'b0;
    defparam \d1.mins_stored_0_sqmuxa_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \d1.mins_stored_0_sqmuxa_LC_10_14_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \d1.mins_stored_0_sqmuxa_LC_10_14_5  (
            .in0(N__11888),
            .in1(N__8796),
            .in2(N__12796),
            .in3(N__8762),
            .lcout(mins_stored_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.secs_0_sqmuxa_ns_LC_10_14_6 .C_ON=1'b0;
    defparam \d1.secs_0_sqmuxa_ns_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \d1.secs_0_sqmuxa_ns_LC_10_14_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \d1.secs_0_sqmuxa_ns_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__10095),
            .in2(_gnd_net_),
            .in3(N__9911),
            .lcout(secs_0_sqmuxa),
            .ltout(secs_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.un1_state_9_LC_10_14_7 .C_ON=1'b0;
    defparam \d1.un1_state_9_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \d1.un1_state_9_LC_10_14_7 .LUT_INIT=16'b0110000001000000;
    LogicCell40 \d1.un1_state_9_LC_10_14_7  (
            .in0(N__11887),
            .in1(N__12789),
            .in2(N__8751),
            .in3(N__9869),
            .lcout(un1_state_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_LC_10_15_1 .C_ON=1'b0;
    defparam \d1.g0_1_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_LC_10_15_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \d1.g0_1_LC_10_15_1  (
            .in0(N__11082),
            .in1(N__9812),
            .in2(N__9012),
            .in3(N__10023),
            .lcout(ten_secs_1_sqmuxa),
            .ltout(ten_secs_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_0_0_1_LC_10_15_2 .C_ON=1'b0;
    defparam \d1.g0_0_0_1_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \d1.g0_0_0_1_LC_10_15_2 .LUT_INIT=16'b1111000100001110;
    LogicCell40 \d1.g0_0_0_1_LC_10_15_2  (
            .in0(N__9000),
            .in1(N__8994),
            .in2(N__8985),
            .in3(N__13631),
            .lcout(),
            .ltout(\d1.g0_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNI7SNV11_LC_10_15_3 .C_ON=1'b0;
    defparam \d1.state_RNI7SNV11_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNI7SNV11_LC_10_15_3 .LUT_INIT=16'b0111100000001111;
    LogicCell40 \d1.state_RNI7SNV11_LC_10_15_3  (
            .in0(N__8982),
            .in1(N__10062),
            .in2(N__8973),
            .in3(N__13543),
            .lcout(),
            .ltout(\d1.un1_mins_4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_1_LC_10_15_4.C_ON=1'b0;
    defparam mins_1_LC_10_15_4.SEQ_MODE=4'b1000;
    defparam mins_1_LC_10_15_4.LUT_INIT=16'b1011100011110000;
    LogicCell40 mins_1_LC_10_15_4 (
            .in0(N__8970),
            .in1(N__11115),
            .in2(N__8964),
            .in3(N__9870),
            .lcout(minsZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14221),
            .ce(),
            .sr(N__11564));
    defparam \d1.count_RNIP9EH_7_LC_10_15_5 .C_ON=1'b0;
    defparam \d1.count_RNIP9EH_7_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIP9EH_7_LC_10_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNIP9EH_7_LC_10_15_5  (
            .in0(N__8961),
            .in1(N__8934),
            .in2(N__8907),
            .in3(N__8877),
            .lcout(\d1.trans_up_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_8_LC_10_16_0 .C_ON=1'b0;
    defparam \d1.g0_8_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \d1.g0_8_LC_10_16_0 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \d1.g0_8_LC_10_16_0  (
            .in0(N__10194),
            .in1(N__8838),
            .in2(N__10826),
            .in3(N__11505),
            .lcout(\d1.un1_mins_1_sqmuxa_0 ),
            .ltout(\d1.un1_mins_1_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNID20IK_3_LC_10_16_1 .C_ON=1'b0;
    defparam \d1.count_RNID20IK_3_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNID20IK_3_LC_10_16_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \d1.count_RNID20IK_3_LC_10_16_1  (
            .in0(N__10911),
            .in1(N__9198),
            .in2(N__8832),
            .in3(N__10163),
            .lcout(),
            .ltout(\d1.un1_mins_3_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI7SNV11_3_LC_10_16_2 .C_ON=1'b0;
    defparam \d1.count_RNI7SNV11_3_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI7SNV11_3_LC_10_16_2 .LUT_INIT=16'b0101000100001000;
    LogicCell40 \d1.count_RNI7SNV11_3_LC_10_16_2  (
            .in0(N__13632),
            .in1(N__13511),
            .in2(N__8829),
            .in3(N__8826),
            .lcout(),
            .ltout(\d1.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_2_LC_10_16_3.C_ON=1'b0;
    defparam mins_2_LC_10_16_3.SEQ_MODE=4'b1000;
    defparam mins_2_LC_10_16_3.LUT_INIT=16'b0011110010101010;
    LogicCell40 mins_2_LC_10_16_3 (
            .in0(N__8820),
            .in1(N__13772),
            .in2(N__8811),
            .in3(N__10892),
            .lcout(minsZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14216),
            .ce(),
            .sr(N__11551));
    defparam \d1.count_RNI0GQ42_7_LC_10_16_4 .C_ON=1'b0;
    defparam \d1.count_RNI0GQ42_7_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI0GQ42_7_LC_10_16_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \d1.count_RNI0GQ42_7_LC_10_16_4  (
            .in0(N__9213),
            .in1(N__10041),
            .in2(N__9207),
            .in3(N__9152),
            .lcout(\d1.g1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIH6847_16_LC_10_17_0 .C_ON=1'b0;
    defparam \d1.count_RNIH6847_16_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIH6847_16_LC_10_17_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \d1.count_RNIH6847_16_LC_10_17_0  (
            .in0(N__9192),
            .in1(N__9180),
            .in2(N__11520),
            .in3(N__10153),
            .lcout(\d1.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI1SGU2_3_LC_10_17_1 .C_ON=1'b0;
    defparam \d1.count_RNI1SGU2_3_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI1SGU2_3_LC_10_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.count_RNI1SGU2_3_LC_10_17_1  (
            .in0(N__9171),
            .in1(N__10946),
            .in2(N__9153),
            .in3(N__9119),
            .lcout(\d1.trans_up_1_0 ),
            .ltout(\d1.trans_up_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNISBML3_LC_10_17_2 .C_ON=1'b0;
    defparam \d1.state_RNISBML3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNISBML3_LC_10_17_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \d1.state_RNISBML3_LC_10_17_2  (
            .in0(N__9080),
            .in1(N__12785),
            .in2(N__9108),
            .in3(N__11904),
            .lcout(\d1.g0_2_0_o2_2 ),
            .ltout(\d1.g0_2_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIA71EK_LC_10_17_3 .C_ON=1'b0;
    defparam \d1.state_RNIA71EK_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIA71EK_LC_10_17_3 .LUT_INIT=16'b1100100000110111;
    LogicCell40 \d1.state_RNIA71EK_LC_10_17_3  (
            .in0(N__10154),
            .in1(N__10061),
            .in2(N__9105),
            .in3(N__13503),
            .lcout(),
            .ltout(\d1.N_19_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_0_LC_10_17_4.C_ON=1'b0;
    defparam mins_0_LC_10_17_4.SEQ_MODE=4'b1000;
    defparam mins_0_LC_10_17_4.LUT_INIT=16'b1111110011101110;
    LogicCell40 mins_0_LC_10_17_4 (
            .in0(N__9102),
            .in1(N__9090),
            .in2(N__9084),
            .in3(N__10897),
            .lcout(minsZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14212),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_2_0_a4_2_LC_10_17_6 .C_ON=1'b0;
    defparam \d1.g0_2_0_a4_2_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \d1.g0_2_0_a4_2_LC_10_17_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \d1.g0_2_0_a4_2_LC_10_17_6  (
            .in0(N__13765),
            .in1(N__13651),
            .in2(N__13535),
            .in3(N__13892),
            .lcout(\d1.g0_2_0_a4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNI4LMC_LC_10_17_7 .C_ON=1'b0;
    defparam \d1.state_RNI4LMC_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNI4LMC_LC_10_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.state_RNI4LMC_LC_10_17_7  (
            .in0(N__13650),
            .in1(N__13499),
            .in2(N__9081),
            .in3(N__13764),
            .lcout(\d1.g2_i_a5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_RNIP8VS_LC_10_18_0 .C_ON=1'b0;
    defparam \d2.sync_1_RNIP8VS_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \d2.sync_1_RNIP8VS_LC_10_18_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \d2.sync_1_RNIP8VS_LC_10_18_0  (
            .in0(N__12246),
            .in1(N__12017),
            .in2(N__11958),
            .in3(N__11752),
            .lcout(\d2.g0_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_6_LC_10_18_1 .C_ON=1'b0;
    defparam \d1.g2_6_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \d1.g2_6_LC_10_18_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \d1.g2_6_LC_10_18_1  (
            .in0(N__11751),
            .in1(N__11945),
            .in2(N__12032),
            .in3(N__12245),
            .lcout(\d1.g2_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNI1DIH_13_LC_10_18_2 .C_ON=1'b0;
    defparam \d2.count_RNI1DIH_13_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNI1DIH_13_LC_10_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNI1DIH_13_LC_10_18_2  (
            .in0(N__11427),
            .in1(N__12151),
            .in2(N__12177),
            .in3(N__11479),
            .lcout(),
            .ltout(\d2.g0_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIJ0PB1_8_LC_10_18_3 .C_ON=1'b0;
    defparam \d2.count_RNIJ0PB1_8_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIJ0PB1_8_LC_10_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNIJ0PB1_8_LC_10_18_3  (
            .in0(N__11165),
            .in1(N__11306),
            .in2(N__9249),
            .in3(N__11221),
            .lcout(),
            .ltout(\d2.g0_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIK9TB3_10_LC_10_18_4 .C_ON=1'b0;
    defparam \d2.count_RNIK9TB3_10_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIK9TB3_10_LC_10_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNIK9TB3_10_LC_10_18_4  (
            .in0(N__12258),
            .in1(N__9246),
            .in2(N__9240),
            .in3(N__9228),
            .lcout(s_dn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_LC_10_18_5 .C_ON=1'b0;
    defparam \d2.state_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \d2.state_LC_10_18_5 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \d2.state_LC_10_18_5  (
            .in0(N__12018),
            .in1(N__11388),
            .in2(N__9222),
            .in3(N__11949),
            .lcout(d2_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14208),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNI3QT21_4_LC_10_18_6 .C_ON=1'b0;
    defparam \d2.count_RNI3QT21_4_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNI3QT21_4_LC_10_18_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d2.count_RNI3QT21_4_LC_10_18_6  (
            .in0(N__11426),
            .in1(N__11480),
            .in2(N__11230),
            .in3(N__11164),
            .lcout(d2_trans_up_1_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_4_LC_10_18_7 .C_ON=1'b0;
    defparam \d1.g2_4_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_4_LC_10_18_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_4_LC_10_18_7  (
            .in0(N__11478),
            .in1(N__11608),
            .in2(N__11761),
            .in3(N__11425),
            .lcout(\d1.g2_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIS7IH_11_LC_10_19_2 .C_ON=1'b0;
    defparam \d2.count_RNIS7IH_11_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIS7IH_11_LC_10_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNIS7IH_11_LC_10_19_2  (
            .in0(N__12135),
            .in1(N__11680),
            .in2(N__12198),
            .in3(N__11620),
            .lcout(\d2.g0_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.state_RNO_0_LC_10_19_3 .C_ON=1'b0;
    defparam \d2.state_RNO_0_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \d2.state_RNO_0_LC_10_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.state_RNO_0_LC_10_19_3  (
            .in0(N__11621),
            .in1(N__12337),
            .in2(N__11697),
            .in3(N__12248),
            .lcout(\d2.trans_up_1_14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_7_LC_10_19_4 .C_ON=1'b0;
    defparam \d1.g2_7_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \d1.g2_7_LC_10_19_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_7_LC_10_19_4  (
            .in0(N__11217),
            .in1(N__11163),
            .in2(N__12348),
            .in3(N__12242),
            .lcout(),
            .ltout(\d1.g2Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_0_3_LC_10_19_5 .C_ON=1'b0;
    defparam \d1.g2_i_a5_0_3_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_0_3_LC_10_19_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \d1.g2_i_a5_0_3_LC_10_19_5  (
            .in0(N__12025),
            .in1(_gnd_net_),
            .in2(N__9372),
            .in3(N__12790),
            .lcout(\d1.g2_i_a5_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_0_a4_7_LC_10_19_6 .C_ON=1'b0;
    defparam \d1.g0_1_0_a4_7_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_0_a4_7_LC_10_19_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \d1.g0_1_0_a4_7_LC_10_19_6  (
            .in0(N__11335),
            .in1(N__13781),
            .in2(N__13546),
            .in3(N__11759),
            .lcout(),
            .ltout(\d1.g0_1_0_a4Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_0_a4_LC_10_19_7 .C_ON=1'b0;
    defparam \d1.g0_1_0_a4_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_0_a4_LC_10_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d1.g0_1_0_a4_LC_10_19_7  (
            .in0(N__11775),
            .in1(N__12113),
            .in2(N__9369),
            .in3(N__11286),
            .lcout(mins_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.un3_count_cry_1_c_LC_11_11_0 .C_ON=1'b1;
    defparam \d4.un3_count_cry_1_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \d4.un3_count_cry_1_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d4.un3_count_cry_1_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__9360),
            .in2(N__9339),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\d4.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d4.count_2_LC_11_11_1 .C_ON=1'b1;
    defparam \d4.count_2_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \d4.count_2_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_2_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__9315),
            .in2(_gnd_net_),
            .in3(N__9303),
            .lcout(\d4.countZ0Z_2 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_1 ),
            .carryout(\d4.un3_count_cry_2 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_3_LC_11_11_2 .C_ON=1'b1;
    defparam \d4.count_3_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \d4.count_3_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_3_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__9300),
            .in2(_gnd_net_),
            .in3(N__9288),
            .lcout(\d4.countZ0Z_3 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_2 ),
            .carryout(\d4.un3_count_cry_3 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_4_LC_11_11_3 .C_ON=1'b1;
    defparam \d4.count_4_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \d4.count_4_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_4_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__9285),
            .in2(_gnd_net_),
            .in3(N__9273),
            .lcout(\d4.countZ0Z_4 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_3 ),
            .carryout(\d4.un3_count_cry_4 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_5_LC_11_11_4 .C_ON=1'b1;
    defparam \d4.count_5_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \d4.count_5_LC_11_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_5_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__9270),
            .in2(_gnd_net_),
            .in3(N__9504),
            .lcout(\d4.countZ0Z_5 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_4 ),
            .carryout(\d4.un3_count_cry_5 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_6_LC_11_11_5 .C_ON=1'b1;
    defparam \d4.count_6_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \d4.count_6_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_6_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__9500),
            .in2(_gnd_net_),
            .in3(N__9486),
            .lcout(\d4.countZ0Z_6 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_5 ),
            .carryout(\d4.un3_count_cry_6 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_7_LC_11_11_6 .C_ON=1'b1;
    defparam \d4.count_7_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \d4.count_7_LC_11_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_7_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__9483),
            .in2(_gnd_net_),
            .in3(N__9471),
            .lcout(\d4.countZ0Z_7 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_6 ),
            .carryout(\d4.un3_count_cry_7 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_8_LC_11_11_7 .C_ON=1'b1;
    defparam \d4.count_8_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \d4.count_8_LC_11_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_8_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__9468),
            .in2(_gnd_net_),
            .in3(N__9456),
            .lcout(\d4.countZ0Z_8 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_7 ),
            .carryout(\d4.un3_count_cry_8 ),
            .clk(N__14241),
            .ce(),
            .sr(N__9620));
    defparam \d4.count_9_LC_11_12_0 .C_ON=1'b1;
    defparam \d4.count_9_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \d4.count_9_LC_11_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_9_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__9453),
            .in2(_gnd_net_),
            .in3(N__9441),
            .lcout(\d4.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\d4.un3_count_cry_9 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_10_LC_11_12_1 .C_ON=1'b1;
    defparam \d4.count_10_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \d4.count_10_LC_11_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_10_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__9437),
            .in2(_gnd_net_),
            .in3(N__9423),
            .lcout(\d4.countZ0Z_10 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_9 ),
            .carryout(\d4.un3_count_cry_10 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_11_LC_11_12_2 .C_ON=1'b1;
    defparam \d4.count_11_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \d4.count_11_LC_11_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_11_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__9420),
            .in2(_gnd_net_),
            .in3(N__9408),
            .lcout(\d4.countZ0Z_11 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_10 ),
            .carryout(\d4.un3_count_cry_11 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_12_LC_11_12_3 .C_ON=1'b1;
    defparam \d4.count_12_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \d4.count_12_LC_11_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_12_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__9404),
            .in2(_gnd_net_),
            .in3(N__9390),
            .lcout(\d4.countZ0Z_12 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_11 ),
            .carryout(\d4.un3_count_cry_12 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_13_LC_11_12_4 .C_ON=1'b1;
    defparam \d4.count_13_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \d4.count_13_LC_11_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_13_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__9387),
            .in2(_gnd_net_),
            .in3(N__9375),
            .lcout(\d4.countZ0Z_13 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_12 ),
            .carryout(\d4.un3_count_cry_13 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_14_LC_11_12_5 .C_ON=1'b1;
    defparam \d4.count_14_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \d4.count_14_LC_11_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_14_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__9671),
            .in2(_gnd_net_),
            .in3(N__9657),
            .lcout(\d4.countZ0Z_14 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_13 ),
            .carryout(\d4.un3_count_cry_14 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_15_LC_11_12_6 .C_ON=1'b1;
    defparam \d4.count_15_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \d4.count_15_LC_11_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d4.count_15_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__9654),
            .in2(_gnd_net_),
            .in3(N__9642),
            .lcout(\d4.countZ0Z_15 ),
            .ltout(),
            .carryin(\d4.un3_count_cry_14 ),
            .carryout(\d4.un3_count_cry_15 ),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d4.count_16_LC_11_12_7 .C_ON=1'b0;
    defparam \d4.count_16_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \d4.count_16_LC_11_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d4.count_16_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__9635),
            .in2(_gnd_net_),
            .in3(N__9639),
            .lcout(\d4.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14236),
            .ce(),
            .sr(N__9621));
    defparam \d3.un3_count_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \d3.un3_count_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \d3.un3_count_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d3.un3_count_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__9606),
            .in2(N__9588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\d3.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_2_LC_11_13_1 .C_ON=1'b1;
    defparam \d3.count_2_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \d3.count_2_LC_11_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_2_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__9567),
            .in2(_gnd_net_),
            .in3(N__9555),
            .lcout(\d3.countZ0Z_2 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_1 ),
            .carryout(\d3.un3_count_cry_2 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_3_LC_11_13_2 .C_ON=1'b1;
    defparam \d3.count_3_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \d3.count_3_LC_11_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_3_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__9552),
            .in2(_gnd_net_),
            .in3(N__9540),
            .lcout(\d3.countZ0Z_3 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_2 ),
            .carryout(\d3.un3_count_cry_3 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_4_LC_11_13_3 .C_ON=1'b1;
    defparam \d3.count_4_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \d3.count_4_LC_11_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_4_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__9537),
            .in2(_gnd_net_),
            .in3(N__9525),
            .lcout(\d3.countZ0Z_4 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_3 ),
            .carryout(\d3.un3_count_cry_4 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_5_LC_11_13_4 .C_ON=1'b1;
    defparam \d3.count_5_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \d3.count_5_LC_11_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_5_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__9521),
            .in2(_gnd_net_),
            .in3(N__9507),
            .lcout(\d3.countZ0Z_5 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_4 ),
            .carryout(\d3.un3_count_cry_5 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_6_LC_11_13_5 .C_ON=1'b1;
    defparam \d3.count_6_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \d3.count_6_LC_11_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_6_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__9801),
            .in2(_gnd_net_),
            .in3(N__9789),
            .lcout(\d3.countZ0Z_6 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_5 ),
            .carryout(\d3.un3_count_cry_6 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_7_LC_11_13_6 .C_ON=1'b1;
    defparam \d3.count_7_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \d3.count_7_LC_11_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_7_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__9786),
            .in2(_gnd_net_),
            .in3(N__9774),
            .lcout(\d3.countZ0Z_7 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_6 ),
            .carryout(\d3.un3_count_cry_7 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_8_LC_11_13_7 .C_ON=1'b1;
    defparam \d3.count_8_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \d3.count_8_LC_11_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_8_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__9771),
            .in2(_gnd_net_),
            .in3(N__9759),
            .lcout(\d3.countZ0Z_8 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_7 ),
            .carryout(\d3.un3_count_cry_8 ),
            .clk(N__14228),
            .ce(),
            .sr(N__9959));
    defparam \d3.count_9_LC_11_14_0 .C_ON=1'b1;
    defparam \d3.count_9_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \d3.count_9_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_9_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__9755),
            .in2(_gnd_net_),
            .in3(N__9741),
            .lcout(\d3.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\d3.un3_count_cry_9 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_10_LC_11_14_1 .C_ON=1'b1;
    defparam \d3.count_10_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \d3.count_10_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_10_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__9737),
            .in2(_gnd_net_),
            .in3(N__9723),
            .lcout(\d3.countZ0Z_10 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_9 ),
            .carryout(\d3.un3_count_cry_10 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_11_LC_11_14_2 .C_ON=1'b1;
    defparam \d3.count_11_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \d3.count_11_LC_11_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_11_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__9716),
            .in2(_gnd_net_),
            .in3(N__9702),
            .lcout(\d3.countZ0Z_11 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_10 ),
            .carryout(\d3.un3_count_cry_11 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_12_LC_11_14_3 .C_ON=1'b1;
    defparam \d3.count_12_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \d3.count_12_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_12_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__9695),
            .in2(_gnd_net_),
            .in3(N__9681),
            .lcout(\d3.countZ0Z_12 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_11 ),
            .carryout(\d3.un3_count_cry_12 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_13_LC_11_14_4 .C_ON=1'b1;
    defparam \d3.count_13_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \d3.count_13_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_13_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__9836),
            .in2(_gnd_net_),
            .in3(N__9678),
            .lcout(\d3.countZ0Z_13 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_12 ),
            .carryout(\d3.un3_count_cry_13 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_14_LC_11_14_5 .C_ON=1'b1;
    defparam \d3.count_14_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \d3.count_14_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_14_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__10632),
            .in2(_gnd_net_),
            .in3(N__9675),
            .lcout(\d3.countZ0Z_14 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_13 ),
            .carryout(\d3.un3_count_cry_14 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_15_LC_11_14_6 .C_ON=1'b1;
    defparam \d3.count_15_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \d3.count_15_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d3.count_15_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__10650),
            .in2(_gnd_net_),
            .in3(N__9966),
            .lcout(\d3.countZ0Z_15 ),
            .ltout(),
            .carryin(\d3.un3_count_cry_14 ),
            .carryout(\d3.un3_count_cry_15 ),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d3.count_16_LC_11_14_7 .C_ON=1'b0;
    defparam \d3.count_16_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \d3.count_16_LC_11_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d3.count_16_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__10668),
            .in2(_gnd_net_),
            .in3(N__9963),
            .lcout(\d3.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14222),
            .ce(),
            .sr(N__9960));
    defparam \d1.un1_state_7_LC_11_15_0 .C_ON=1'b0;
    defparam \d1.un1_state_7_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \d1.un1_state_7_LC_11_15_0 .LUT_INIT=16'b0011100000000000;
    LogicCell40 \d1.un1_state_7_LC_11_15_0  (
            .in0(N__9868),
            .in1(N__11891),
            .in2(N__12801),
            .in3(N__9945),
            .lcout(un1_state_7_0),
            .ltout(un1_state_7_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_1_LC_11_15_1.C_ON=1'b0;
    defparam secs_1_LC_11_15_1.SEQ_MODE=4'b1000;
    defparam secs_1_LC_11_15_1.LUT_INIT=16'b1001101000000000;
    LogicCell40 secs_1_LC_11_15_1 (
            .in0(N__10442),
            .in1(N__10351),
            .in2(N__9882),
            .in3(N__9876),
            .lcout(secsZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14217),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.un1_alarm_on_0_sqmuxa_0_i_LC_11_15_2 .C_ON=1'b0;
    defparam \d1.un1_alarm_on_0_sqmuxa_0_i_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \d1.un1_alarm_on_0_sqmuxa_0_i_LC_11_15_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \d1.un1_alarm_on_0_sqmuxa_0_i_LC_11_15_2  (
            .in0(N__12795),
            .in1(N__9866),
            .in2(_gnd_net_),
            .in3(N__11889),
            .lcout(un1_alarm_on_0_sqmuxa_0_i),
            .ltout(un1_alarm_on_0_sqmuxa_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_RNO_0_1_LC_11_15_3.C_ON=1'b0;
    defparam secs_RNO_0_1_LC_11_15_3.SEQ_MODE=4'b0000;
    defparam secs_RNO_0_1_LC_11_15_3.LUT_INIT=16'b0000001100001111;
    LogicCell40 secs_RNO_0_1_LC_11_15_3 (
            .in0(_gnd_net_),
            .in1(N__10534),
            .in2(N__9879),
            .in3(N__10025),
            .lcout(N_120_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_0_sqmuxa_1_LC_11_15_4 .C_ON=1'b0;
    defparam \d1.state_0_sqmuxa_1_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \d1.state_0_sqmuxa_1_LC_11_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \d1.state_0_sqmuxa_1_LC_11_15_4  (
            .in0(N__13542),
            .in1(N__13866),
            .in2(N__13634),
            .in3(N__13776),
            .lcout(\d1.state_0_sqmuxaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_2_LC_11_15_5 .C_ON=1'b0;
    defparam \d1.g0_2_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \d1.g0_2_LC_11_15_5 .LUT_INIT=16'b1001100111111111;
    LogicCell40 \d1.g0_2_LC_11_15_5  (
            .in0(N__11890),
            .in1(N__12791),
            .in2(_gnd_net_),
            .in3(N__9867),
            .lcout(un1_alarm_on_0_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.state_RNI607I1_LC_11_15_6 .C_ON=1'b0;
    defparam \d3.state_RNI607I1_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \d3.state_RNI607I1_LC_11_15_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \d3.state_RNI607I1_LC_11_15_6  (
            .in0(N__12567),
            .in1(N__9832),
            .in2(N__12617),
            .in3(N__10614),
            .lcout(d3_g0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.secs_0_sqmuxa_x1_LC_11_15_7 .C_ON=1'b0;
    defparam \d1.secs_0_sqmuxa_x1_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \d1.secs_0_sqmuxa_x1_LC_11_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \d1.secs_0_sqmuxa_x1_LC_11_15_7  (
            .in0(N__10469),
            .in1(N__10435),
            .in2(N__10399),
            .in3(N__10350),
            .lcout(\d1.secs_0_sqmuxa_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.mins_16_1_3_LC_11_16_0 .C_ON=1'b0;
    defparam \d1.mins_16_1_3_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \d1.mins_16_1_3_LC_11_16_0 .LUT_INIT=16'b0100011110001011;
    LogicCell40 \d1.mins_16_1_3_LC_11_16_0  (
            .in0(N__13849),
            .in1(N__10878),
            .in2(N__10086),
            .in3(N__10060),
            .lcout(\d1.mins_16_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_0_LC_11_16_1.C_ON=1'b0;
    defparam secs_0_LC_11_16_1.SEQ_MODE=4'b1000;
    defparam secs_0_LC_11_16_1.LUT_INIT=16'b0000000001100110;
    LogicCell40 secs_0_LC_11_16_1 (
            .in0(N__10358),
            .in1(N__9999),
            .in2(_gnd_net_),
            .in3(N__9976),
            .lcout(secsZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14213),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIC9AJK_16_LC_11_16_2 .C_ON=1'b0;
    defparam \d1.count_RNIC9AJK_16_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIC9AJK_16_LC_11_16_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \d1.count_RNIC9AJK_16_LC_11_16_2  (
            .in0(N__13510),
            .in1(N__10068),
            .in2(N__12522),
            .in3(N__10059),
            .lcout(\d1.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_10_LC_11_16_3 .C_ON=1'b0;
    defparam \d1.g0_10_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \d1.g0_10_LC_11_16_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \d1.g0_10_LC_11_16_3  (
            .in0(N__13487),
            .in1(N__13848),
            .in2(N__13680),
            .in3(N__13755),
            .lcout(\d1.g0_0_0_a4_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_RNO_0_2_LC_11_16_4.C_ON=1'b0;
    defparam secs_RNO_0_2_LC_11_16_4.SEQ_MODE=4'b0000;
    defparam secs_RNO_0_2_LC_11_16_4.LUT_INIT=16'b1010101010011010;
    LogicCell40 secs_RNO_0_2_LC_11_16_4 (
            .in0(N__10473),
            .in1(N__10440),
            .in2(N__10001),
            .in3(N__10356),
            .lcout(),
            .ltout(secs_RNO_0Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_2_LC_11_16_5.C_ON=1'b0;
    defparam secs_2_LC_11_16_5.SEQ_MODE=4'b1000;
    defparam secs_2_LC_11_16_5.LUT_INIT=16'b0001000000110000;
    LogicCell40 secs_2_LC_11_16_5 (
            .in0(N__10550),
            .in1(N__9978),
            .in2(N__10032),
            .in3(N__10029),
            .lcout(secsZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14213),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_RNO_0_3_LC_11_16_6.C_ON=1'b0;
    defparam secs_RNO_0_3_LC_11_16_6.SEQ_MODE=4'b0000;
    defparam secs_RNO_0_3_LC_11_16_6.LUT_INIT=16'b1111000011100000;
    LogicCell40 secs_RNO_0_3_LC_11_16_6 (
            .in0(N__10474),
            .in1(N__10441),
            .in2(N__10002),
            .in3(N__10357),
            .lcout(),
            .ltout(un1_secs_c3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_3_LC_11_16_7.C_ON=1'b0;
    defparam secs_3_LC_11_16_7.SEQ_MODE=4'b1000;
    defparam secs_3_LC_11_16_7.LUT_INIT=16'b0000000010010110;
    LogicCell40 secs_3_LC_11_16_7 (
            .in0(N__10398),
            .in1(N__10000),
            .in2(N__9981),
            .in3(N__9977),
            .lcout(secsZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14213),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIGDI57_LC_11_17_0 .C_ON=1'b0;
    defparam \d1.state_RNIGDI57_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIGDI57_LC_11_17_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \d1.state_RNIGDI57_LC_11_17_0  (
            .in0(N__10217),
            .in1(N__10101),
            .in2(N__10206),
            .in3(N__11370),
            .lcout(\d1.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_9_LC_11_17_1 .C_ON=1'b0;
    defparam \d1.g0_9_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \d1.g0_9_LC_11_17_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \d1.g0_9_LC_11_17_1  (
            .in0(N__13748),
            .in1(N__13488),
            .in2(N__13681),
            .in3(N__13850),
            .lcout(\d1.mins27_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_0_1_LC_11_17_2 .C_ON=1'b0;
    defparam \d1.g0_0_1_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \d1.g0_0_1_LC_11_17_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \d1.g0_0_1_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__13841),
            .in2(_gnd_net_),
            .in3(N__13747),
            .lcout(),
            .ltout(\d1.g0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_10_LC_11_17_3 .C_ON=1'b0;
    defparam \d1.g2_10_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \d1.g2_10_LC_11_17_3 .LUT_INIT=16'b0100000011111111;
    LogicCell40 \d1.g2_10_LC_11_17_3  (
            .in0(N__13670),
            .in1(N__13489),
            .in2(N__10197),
            .in3(N__11269),
            .lcout(\d1.g2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIINS67_0_LC_11_17_4 .C_ON=1'b0;
    defparam \d1.state_RNIINS67_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIINS67_0_LC_11_17_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \d1.state_RNIINS67_0_LC_11_17_4  (
            .in0(N__10187),
            .in1(N__10162),
            .in2(_gnd_net_),
            .in3(N__10125),
            .lcout(\d1.mins_2_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_0_6_LC_11_17_5 .C_ON=1'b0;
    defparam \d1.g2_i_a5_0_6_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_0_6_LC_11_17_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \d1.g2_i_a5_0_6_LC_11_17_5  (
            .in0(N__11696),
            .in1(N__10113),
            .in2(N__11985),
            .in3(N__11900),
            .lcout(),
            .ltout(\d1.g2_i_a5_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_0_LC_11_17_6 .C_ON=1'b0;
    defparam \d1.g2_i_0_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_0_LC_11_17_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \d1.g2_i_0_LC_11_17_6  (
            .in0(N__11349),
            .in1(N__11313),
            .in2(N__10104),
            .in3(N__12054),
            .lcout(\d1.g2_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_2_LC_11_17_7 .C_ON=1'b0;
    defparam \d1.g2_i_a5_2_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_2_LC_11_17_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \d1.g2_i_a5_2_LC_11_17_7  (
            .in0(N__12784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11899),
            .lcout(\d1.g2_i_a5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.un3_count_cry_1_c_LC_11_18_0 .C_ON=1'b1;
    defparam \d2.un3_count_cry_1_c_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \d2.un3_count_cry_1_c_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \d2.un3_count_cry_1_c_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__11448),
            .in2(N__11643),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\d2.un3_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_2_LC_11_18_1 .C_ON=1'b1;
    defparam \d2.count_2_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \d2.count_2_LC_11_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_2_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__11694),
            .in2(_gnd_net_),
            .in3(N__10248),
            .lcout(d2_count_2),
            .ltout(),
            .carryin(\d2.un3_count_cry_1 ),
            .carryout(\d2.un3_count_cry_2 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_3_LC_11_18_2 .C_ON=1'b1;
    defparam \d2.count_3_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \d2.count_3_LC_11_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_3_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__12247),
            .in2(_gnd_net_),
            .in3(N__10245),
            .lcout(d2_count_3),
            .ltout(),
            .carryin(\d2.un3_count_cry_2 ),
            .carryout(\d2.un3_count_cry_3 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_4_LC_11_18_3 .C_ON=1'b1;
    defparam \d2.count_4_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \d2.count_4_LC_11_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_4_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__11488),
            .in2(_gnd_net_),
            .in3(N__10242),
            .lcout(d2_count_4),
            .ltout(),
            .carryin(\d2.un3_count_cry_3 ),
            .carryout(\d2.un3_count_cry_4 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_5_LC_11_18_4 .C_ON=1'b1;
    defparam \d2.count_5_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \d2.count_5_LC_11_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_5_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__11172),
            .in2(_gnd_net_),
            .in3(N__10239),
            .lcout(d2_count_5),
            .ltout(),
            .carryin(\d2.un3_count_cry_4 ),
            .carryout(\d2.un3_count_cry_5 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_6_LC_11_18_5 .C_ON=1'b1;
    defparam \d2.count_6_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \d2.count_6_LC_11_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_6_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__11228),
            .in2(_gnd_net_),
            .in3(N__10236),
            .lcout(d2_count_6),
            .ltout(),
            .carryin(\d2.un3_count_cry_5 ),
            .carryout(\d2.un3_count_cry_6 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_7_LC_11_18_6 .C_ON=1'b1;
    defparam \d2.count_7_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \d2.count_7_LC_11_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_7_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__12273),
            .in2(_gnd_net_),
            .in3(N__10233),
            .lcout(\d2.countZ0Z_7 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_6 ),
            .carryout(\d2.un3_count_cry_7 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_8_LC_11_18_7 .C_ON=1'b1;
    defparam \d2.count_8_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_8_LC_11_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_8_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__11307),
            .in2(_gnd_net_),
            .in3(N__10230),
            .lcout(\d2.countZ0Z_8 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_7 ),
            .carryout(\d2.un3_count_cry_8 ),
            .clk(N__14205),
            .ce(),
            .sr(N__10289));
    defparam \d2.count_9_LC_11_19_0 .C_ON=1'b1;
    defparam \d2.count_9_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \d2.count_9_LC_11_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_9_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__12372),
            .in2(_gnd_net_),
            .in3(N__10227),
            .lcout(\d2.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\d2.un3_count_cry_9 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_10_LC_11_19_1 .C_ON=1'b1;
    defparam \d2.count_10_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \d2.count_10_LC_11_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_10_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__12292),
            .in2(_gnd_net_),
            .in3(N__10224),
            .lcout(\d2.countZ0Z_10 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_9 ),
            .carryout(\d2.un3_count_cry_10 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_11_LC_11_19_2 .C_ON=1'b1;
    defparam \d2.count_11_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \d2.count_11_LC_11_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_11_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__12134),
            .in2(_gnd_net_),
            .in3(N__10308),
            .lcout(\d2.countZ0Z_11 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_10 ),
            .carryout(\d2.un3_count_cry_11 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_12_LC_11_19_3 .C_ON=1'b1;
    defparam \d2.count_12_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \d2.count_12_LC_11_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_12_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__12197),
            .in2(_gnd_net_),
            .in3(N__10305),
            .lcout(\d2.countZ0Z_12 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_11 ),
            .carryout(\d2.un3_count_cry_12 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_13_LC_11_19_4 .C_ON=1'b1;
    defparam \d2.count_13_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \d2.count_13_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_13_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__12176),
            .in2(_gnd_net_),
            .in3(N__10302),
            .lcout(\d2.countZ0Z_13 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_12 ),
            .carryout(\d2.un3_count_cry_13 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_14_LC_11_19_5 .C_ON=1'b1;
    defparam \d2.count_14_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \d2.count_14_LC_11_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_14_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__12155),
            .in2(_gnd_net_),
            .in3(N__10299),
            .lcout(\d2.countZ0Z_14 ),
            .ltout(),
            .carryin(\d2.un3_count_cry_13 ),
            .carryout(\d2.un3_count_cry_14 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_15_LC_11_19_6 .C_ON=1'b1;
    defparam \d2.count_15_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \d2.count_15_LC_11_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \d2.count_15_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__11760),
            .in2(_gnd_net_),
            .in3(N__10296),
            .lcout(d2_count_15),
            .ltout(),
            .carryin(\d2.un3_count_cry_14 ),
            .carryout(\d2.un3_count_cry_15 ),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam \d2.count_16_LC_11_19_7 .C_ON=1'b0;
    defparam \d2.count_16_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \d2.count_16_LC_11_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \d2.count_16_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__12341),
            .in2(_gnd_net_),
            .in3(N__10293),
            .lcout(d2_count_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14204),
            .ce(),
            .sr(N__10288));
    defparam state_e_1_LC_12_12_0.C_ON=1'b0;
    defparam state_e_1_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam state_e_1_LC_12_12_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 state_e_1_LC_12_12_0 (
            .in0(N__10731),
            .in1(N__10323),
            .in2(_gnd_net_),
            .in3(N__10549),
            .lcout(stateZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14223),
            .ce(N__10275),
            .sr(_gnd_net_));
    defparam state_sbtinv_1_LC_12_13_5.C_ON=1'b0;
    defparam state_sbtinv_1_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam state_sbtinv_1_LC_12_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 state_sbtinv_1_LC_12_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10254),
            .lcout(un1_state_0_sqmuxa_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.un1_state_0_sqmuxa_1_LC_12_13_6 .C_ON=1'b0;
    defparam \d1.un1_state_0_sqmuxa_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \d1.un1_state_0_sqmuxa_1_LC_12_13_6 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \d1.un1_state_0_sqmuxa_1_LC_12_13_6  (
            .in0(N__10719),
            .in1(N__10263),
            .in2(N__10545),
            .in3(N__10710),
            .lcout(un1_state_0_sqmuxa_1_0),
            .ltout(un1_state_0_sqmuxa_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state_0_LC_12_13_7.C_ON=1'b0;
    defparam state_0_LC_12_13_7.SEQ_MODE=4'b1001;
    defparam state_0_LC_12_13_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 state_0_LC_12_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10782),
            .in3(N__12716),
            .lcout(stateZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14218),
            .ce(),
            .sr(N__10779));
    defparam \d1.state_0_sqmuxa_2_LC_12_14_0 .C_ON=1'b0;
    defparam \d1.state_0_sqmuxa_2_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \d1.state_0_sqmuxa_2_LC_12_14_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \d1.state_0_sqmuxa_2_LC_12_14_0  (
            .in0(N__10608),
            .in1(N__12495),
            .in2(N__10743),
            .in3(N__12450),
            .lcout(\d1.state_0_sqmuxaZ0Z_2 ),
            .ltout(\d1.state_0_sqmuxaZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_0_sqmuxa_LC_12_14_1 .C_ON=1'b0;
    defparam \d1.state_0_sqmuxa_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \d1.state_0_sqmuxa_LC_12_14_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \d1.state_0_sqmuxa_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__10319),
            .in2(N__10722),
            .in3(N__10530),
            .lcout(state_0_sqmuxa),
            .ltout(state_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam alarm_on_LC_12_14_2.C_ON=1'b0;
    defparam alarm_on_LC_12_14_2.SEQ_MODE=4'b1000;
    defparam alarm_on_LC_12_14_2.LUT_INIT=16'b1111000011111100;
    LogicCell40 alarm_on_LC_12_14_2 (
            .in0(_gnd_net_),
            .in1(N__10682),
            .in2(N__10713),
            .in3(N__10709),
            .lcout(alarm_onZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14214),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.count_RNI4GDS_16_LC_12_14_3 .C_ON=1'b0;
    defparam \d3.count_RNI4GDS_16_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \d3.count_RNI4GDS_16_LC_12_14_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \d3.count_RNI4GDS_16_LC_12_14_3  (
            .in0(N__10667),
            .in1(N__10648),
            .in2(_gnd_net_),
            .in3(N__10630),
            .lcout(\d3.count_RNI4GDSZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.un1_state_3_LC_12_14_7 .C_ON=1'b0;
    defparam \d1.un1_state_3_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \d1.un1_state_3_LC_12_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \d1.un1_state_3_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__11860),
            .in2(_gnd_net_),
            .in3(N__12684),
            .lcout(un1_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_0_2_LC_12_15_0 .C_ON=1'b0;
    defparam \d1.g0_0_2_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \d1.g0_0_2_LC_12_15_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \d1.g0_0_2_LC_12_15_0  (
            .in0(N__10599),
            .in1(N__12505),
            .in2(N__10544),
            .in3(N__12451),
            .lcout(\d1.g0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secs_RNIUG5J_3_LC_12_15_3.C_ON=1'b0;
    defparam secs_RNIUG5J_3_LC_12_15_3.SEQ_MODE=4'b0000;
    defparam secs_RNIUG5J_3_LC_12_15_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 secs_RNIUG5J_3_LC_12_15_3 (
            .in0(N__10478),
            .in1(N__10436),
            .in2(N__10400),
            .in3(N__10352),
            .lcout(decrement_time_0_secs9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_3_LC_12_15_4 .C_ON=1'b0;
    defparam \d1.g2_3_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \d1.g2_3_LC_12_15_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_3_LC_12_15_4  (
            .in0(N__11229),
            .in1(N__11173),
            .in2(N__12357),
            .in3(N__12249),
            .lcout(),
            .ltout(\d1.g2_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_1_LC_12_15_5 .C_ON=1'b0;
    defparam \d1.g2_1_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \d1.g2_1_LC_12_15_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \d1.g2_1_LC_12_15_5  (
            .in0(N__12047),
            .in1(N__11981),
            .in2(N__11127),
            .in3(N__11861),
            .lcout(\d1.g2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_13_LC_12_15_6 .C_ON=1'b0;
    defparam \d1.g2_13_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \d1.g2_13_LC_12_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \d1.g2_13_LC_12_15_6  (
            .in0(N__11862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12749),
            .lcout(\d1.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.state_LC_12_15_7 .C_ON=1'b0;
    defparam \d3.state_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \d3.state_LC_12_15_7 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \d3.state_LC_12_15_7  (
            .in0(N__12618),
            .in1(N__12575),
            .in2(N__11106),
            .in3(N__11091),
            .lcout(\d3.stateZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14209),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNI2PCE_1_3_LC_12_16_0 .C_ON=1'b0;
    defparam \d1.count_RNI2PCE_1_3_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNI2PCE_1_3_LC_12_16_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.count_RNI2PCE_1_3_LC_12_16_0  (
            .in0(N__11061),
            .in1(N__11034),
            .in2(N__11007),
            .in3(N__10974),
            .lcout(),
            .ltout(\d1.g1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.count_RNIUT4M1_3_LC_12_16_1 .C_ON=1'b0;
    defparam \d1.count_RNIUT4M1_3_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \d1.count_RNIUT4M1_3_LC_12_16_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \d1.count_RNIUT4M1_3_LC_12_16_1  (
            .in0(N__10950),
            .in1(N__11901),
            .in2(N__10914),
            .in3(N__12748),
            .lcout(\d1.g1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.state_RNIKMMMV_LC_12_16_5 .C_ON=1'b0;
    defparam \d1.state_RNIKMMMV_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \d1.state_RNIKMMMV_LC_12_16_5 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \d1.state_RNIKMMMV_LC_12_16_5  (
            .in0(N__10885),
            .in1(N__10845),
            .in2(N__10839),
            .in3(N__10830),
            .lcout(),
            .ltout(\d1.g3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mins_3_LC_12_16_6.C_ON=1'b0;
    defparam mins_3_LC_12_16_6.SEQ_MODE=4'b1001;
    defparam mins_3_LC_12_16_6.LUT_INIT=16'b0001010000010001;
    LogicCell40 mins_3_LC_12_16_6 (
            .in0(N__10803),
            .in1(N__10797),
            .in2(N__10791),
            .in3(N__10788),
            .lcout(minsZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14206),
            .ce(),
            .sr(N__11568));
    defparam \d1.g0_1_a5_0_11_LC_12_17_0 .C_ON=1'b0;
    defparam \d1.g0_1_a5_0_11_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_a5_0_11_LC_12_17_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \d1.g0_1_a5_0_11_LC_12_17_0  (
            .in0(N__12774),
            .in1(N__13862),
            .in2(N__13548),
            .in3(N__11898),
            .lcout(\d1.g0_1_a5_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_14_LC_12_17_1 .C_ON=1'b0;
    defparam \d1.g2_14_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \d1.g2_14_LC_12_17_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \d1.g2_14_LC_12_17_1  (
            .in0(N__12100),
            .in1(N__12204),
            .in2(N__12797),
            .in3(N__12352),
            .lcout(\d1.g2_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_8_LC_12_17_3 .C_ON=1'b0;
    defparam \d1.g2_8_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \d1.g2_8_LC_12_17_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \d1.g2_8_LC_12_17_3  (
            .in0(N__11484),
            .in1(N__11638),
            .in2(N__11766),
            .in3(N__11447),
            .lcout(\d1.g2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNID7FT1_15_LC_12_17_4 .C_ON=1'b0;
    defparam \d2.count_RNID7FT1_15_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNID7FT1_15_LC_12_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \d2.count_RNID7FT1_15_LC_12_17_4  (
            .in0(N__11343),
            .in1(N__11765),
            .in2(N__12102),
            .in3(N__11270),
            .lcout(\d2.trans_up_1_15 ),
            .ltout(\d2.trans_up_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIK9TB3_1_LC_12_17_5 .C_ON=1'b0;
    defparam \d2.count_RNIK9TB3_1_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIK9TB3_1_LC_12_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNIK9TB3_1_LC_12_17_5  (
            .in0(N__11919),
            .in1(N__11639),
            .in2(N__11373),
            .in3(N__11695),
            .lcout(s_dn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_0_7_LC_12_17_6 .C_ON=1'b0;
    defparam \d1.g2_i_a5_0_7_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_0_7_LC_12_17_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \d1.g2_i_a5_0_7_LC_12_17_6  (
            .in0(N__11364),
            .in1(N__12101),
            .in2(N__11358),
            .in3(N__11271),
            .lcout(\d1.g2_i_a5_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIQ9VS_16_LC_12_18_0 .C_ON=1'b0;
    defparam \d2.count_RNIQ9VS_16_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIQ9VS_16_LC_12_18_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \d2.count_RNIQ9VS_16_LC_12_18_0  (
            .in0(N__12244),
            .in1(N__11973),
            .in2(N__12046),
            .in3(N__12327),
            .lcout(d2_g0_3),
            .ltout(d2_g0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_1_7_LC_12_18_1 .C_ON=1'b0;
    defparam \d1.g2_i_a5_1_7_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_1_7_LC_12_18_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \d1.g2_i_a5_1_7_LC_12_18_1  (
            .in0(N__12096),
            .in1(N__11342),
            .in2(N__11316),
            .in3(N__11272),
            .lcout(\d1.g2_i_a5_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNITE8Q_10_LC_12_18_2 .C_ON=1'b0;
    defparam \d2.count_RNITE8Q_10_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNITE8Q_10_LC_12_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNITE8Q_10_LC_12_18_2  (
            .in0(N__12370),
            .in1(N__11299),
            .in2(N__12293),
            .in3(N__12271),
            .lcout(d2_trans_up_1_15_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNICOIH_10_LC_12_18_4 .C_ON=1'b0;
    defparam \d2.count_RNICOIH_10_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNICOIH_10_LC_12_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNICOIH_10_LC_12_18_4  (
            .in0(N__12371),
            .in1(N__12326),
            .in2(N__12294),
            .in3(N__12272),
            .lcout(\d2.g0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_16_LC_12_18_5 .C_ON=1'b0;
    defparam \d1.g2_16_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \d1.g2_16_LC_12_18_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \d1.g2_16_LC_12_18_5  (
            .in0(N__11972),
            .in1(N__11753),
            .in2(N__12045),
            .in3(N__12243),
            .lcout(\d1.g2_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNI237_11_LC_12_18_6 .C_ON=1'b0;
    defparam \d2.count_RNI237_11_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNI237_11_LC_12_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \d2.count_RNI237_11_LC_12_18_6  (
            .in0(N__12193),
            .in1(N__12175),
            .in2(N__12156),
            .in3(N__12130),
            .lcout(d2_trans_up_1_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_1_6_LC_12_18_7 .C_ON=1'b0;
    defparam \d1.g2_i_a5_1_6_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_1_6_LC_12_18_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \d1.g2_i_a5_1_6_LC_12_18_7  (
            .in0(N__13550),
            .in1(N__12624),
            .in2(N__13682),
            .in3(N__11864),
            .lcout(\d1.g2_i_a5_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.sync_1_RNIMV5K_LC_12_19_1 .C_ON=1'b0;
    defparam \d2.sync_1_RNIMV5K_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \d2.sync_1_RNIMV5K_LC_12_19_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \d2.sync_1_RNIMV5K_LC_12_19_1  (
            .in0(N__12048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11980),
            .lcout(\d2.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_0_a4_4_LC_12_19_4 .C_ON=1'b0;
    defparam \d1.g0_1_0_a4_4_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_0_a4_4_LC_12_19_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \d1.g0_1_0_a4_4_LC_12_19_4  (
            .in0(N__13867),
            .in1(N__11684),
            .in2(N__13679),
            .in3(N__11628),
            .lcout(),
            .ltout(\d1.g0_1_0_a4Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_0_a4_8_LC_12_19_5 .C_ON=1'b0;
    defparam \d1.g0_1_0_a4_8_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_0_a4_8_LC_12_19_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \d1.g0_1_0_a4_8_LC_12_19_5  (
            .in0(N__11918),
            .in1(N__12731),
            .in2(N__11907),
            .in3(N__11863),
            .lcout(\d1.g0_1_0_a4Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d2.count_RNIOJGH_15_LC_12_19_6 .C_ON=1'b0;
    defparam \d2.count_RNIOJGH_15_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \d2.count_RNIOJGH_15_LC_12_19_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \d2.count_RNIOJGH_15_LC_12_19_6  (
            .in0(N__11747),
            .in1(N__11685),
            .in2(_gnd_net_),
            .in3(N__11627),
            .lcout(),
            .ltout(d2_g0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g2_i_a5_1_3_LC_12_19_7 .C_ON=1'b0;
    defparam \d1.g2_i_a5_1_3_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \d1.g2_i_a5_1_3_LC_12_19_7 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \d1.g2_i_a5_1_3_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__12732),
            .in2(N__12627),
            .in3(N__13789),
            .lcout(\d1.g2_i_a5_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_8_LC_13_13_0 .C_ON=1'b0;
    defparam \display2.prescaler_8_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_8_LC_13_13_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display2.prescaler_8_LC_13_13_0  (
            .in0(N__13984),
            .in1(N__13074),
            .in2(N__14043),
            .in3(N__12813),
            .lcout(\display2.prescalerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14229),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNI3D3L_23_LC_13_13_1 .C_ON=1'b0;
    defparam \display2.prescaler_RNI3D3L_23_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNI3D3L_23_LC_13_13_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \display2.prescaler_RNI3D3L_23_LC_13_13_1  (
            .in0(N__12824),
            .in1(N__12848),
            .in2(N__13017),
            .in3(N__12872),
            .lcout(\display2.prescaler8_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_6_LC_13_13_3 .C_ON=1'b0;
    defparam \display2.prescaler_6_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_6_LC_13_13_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \display2.prescaler_6_LC_13_13_3  (
            .in0(N__12837),
            .in1(N__14038),
            .in2(N__13083),
            .in3(N__13983),
            .lcout(\display2.prescalerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14229),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_4_LC_13_13_5 .C_ON=1'b0;
    defparam \display2.prescaler_4_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_4_LC_13_13_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \display2.prescaler_4_LC_13_13_5  (
            .in0(N__12861),
            .in1(N__14037),
            .in2(N__13082),
            .in3(N__13982),
            .lcout(\display2.prescalerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14229),
            .ce(),
            .sr(_gnd_net_));
    defparam \d3.state_RNIOCAC_LC_13_14_2 .C_ON=1'b0;
    defparam \d3.state_RNIOCAC_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \d3.state_RNIOCAC_LC_13_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \d3.state_RNIOCAC_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__12610),
            .in2(_gnd_net_),
            .in3(N__12568),
            .lcout(\d3.idle_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.g0_1_0_0_LC_13_14_7 .C_ON=1'b0;
    defparam \d1.g0_1_0_0_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \d1.g0_1_0_0_LC_13_14_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \d1.g0_1_0_0_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__13675),
            .in2(_gnd_net_),
            .in3(N__13790),
            .lcout(\d1.g0_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.BNC1_LC_13_16_1 .C_ON=1'b0;
    defparam \d1.BNC1_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \d1.BNC1_LC_13_16_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \d1.BNC1_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__12506),
            .in2(_gnd_net_),
            .in3(N__12452),
            .lcout(BNC1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_2_cry_1_c_LC_14_12_0 .C_ON=1'b1;
    defparam \display2.prescaler_2_cry_1_c_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_2_cry_1_c_LC_14_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \display2.prescaler_2_cry_1_c_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__13101),
            .in2(N__13206),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\display2.prescaler_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_2_LC_14_12_1 .C_ON=1'b1;
    defparam \display2.prescaler_2_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_2_LC_14_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_2_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__12918),
            .in2(_gnd_net_),
            .in3(N__12879),
            .lcout(\display2.prescalerZ0Z_2 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_1 ),
            .carryout(\display2.prescaler_2_cry_2 ),
            .clk(N__14242),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_3_LC_14_12_2 .C_ON=1'b1;
    defparam \display2.prescaler_3_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_3_LC_14_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_3_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__12945),
            .in2(_gnd_net_),
            .in3(N__12876),
            .lcout(\display2.prescalerZ0Z_3 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_2 ),
            .carryout(\display2.prescaler_2_cry_3 ),
            .clk(N__14242),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_4_LC_14_12_3 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_4_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_4_LC_14_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_4_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__12873),
            .in2(_gnd_net_),
            .in3(N__12855),
            .lcout(\display2.prescaler_2_4 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_3 ),
            .carryout(\display2.prescaler_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_5_LC_14_12_4 .C_ON=1'b1;
    defparam \display2.prescaler_5_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_5_LC_14_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_5_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__12957),
            .in2(_gnd_net_),
            .in3(N__12852),
            .lcout(\display2.prescalerZ0Z_5 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_4 ),
            .carryout(\display2.prescaler_2_cry_5 ),
            .clk(N__14242),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_6_LC_14_12_5 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_6_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_6_LC_14_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_6_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__12849),
            .in2(_gnd_net_),
            .in3(N__12831),
            .lcout(\display2.prescaler_2_6 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_5 ),
            .carryout(\display2.prescaler_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_7_LC_14_12_6 .C_ON=1'b1;
    defparam \display2.prescaler_7_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_7_LC_14_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_7_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__12932),
            .in2(_gnd_net_),
            .in3(N__12828),
            .lcout(\display2.prescalerZ0Z_7 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_6 ),
            .carryout(\display2.prescaler_2_cry_7 ),
            .clk(N__14242),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_8_LC_14_12_7 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_8_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_8_LC_14_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_8_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__12825),
            .in2(_gnd_net_),
            .in3(N__12807),
            .lcout(\display2.prescaler_2_8 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_7 ),
            .carryout(\display2.prescaler_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_9_LC_14_13_0 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_9_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_9_LC_14_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_9_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__13173),
            .in2(_gnd_net_),
            .in3(N__12804),
            .lcout(\display2.prescaler_2_9 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\display2.prescaler_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_10_LC_14_13_1 .C_ON=1'b1;
    defparam \display2.prescaler_10_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_10_LC_14_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_10_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__13269),
            .in2(_gnd_net_),
            .in3(N__12906),
            .lcout(\display2.prescalerZ0Z_10 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_9 ),
            .carryout(\display2.prescaler_2_cry_10 ),
            .clk(N__14237),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_11_LC_14_13_2 .C_ON=1'b1;
    defparam \display2.prescaler_11_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_11_LC_14_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_11_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__13239),
            .in2(_gnd_net_),
            .in3(N__12903),
            .lcout(\display2.prescalerZ0Z_11 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_10 ),
            .carryout(\display2.prescaler_2_cry_11 ),
            .clk(N__14237),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_12_LC_14_13_3 .C_ON=1'b1;
    defparam \display2.prescaler_12_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_12_LC_14_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_12_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__13283),
            .in2(_gnd_net_),
            .in3(N__12900),
            .lcout(\display2.prescalerZ0Z_12 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_11 ),
            .carryout(\display2.prescaler_2_cry_12 ),
            .clk(N__14237),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_13_LC_14_13_4 .C_ON=1'b1;
    defparam \display2.prescaler_13_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_13_LC_14_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_13_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__13253),
            .in2(_gnd_net_),
            .in3(N__12897),
            .lcout(\display2.prescalerZ0Z_13 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_12 ),
            .carryout(\display2.prescaler_2_cry_13 ),
            .clk(N__14237),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_14_LC_14_13_5 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_14_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_14_LC_14_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_14_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__13155),
            .in2(_gnd_net_),
            .in3(N__12894),
            .lcout(\display2.prescaler_2_14 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_13 ),
            .carryout(\display2.prescaler_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNO_0_15_LC_14_13_6 .C_ON=1'b1;
    defparam \display2.prescaler_RNO_0_15_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNO_0_15_LC_14_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_RNO_0_15_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__13952),
            .in2(_gnd_net_),
            .in3(N__12891),
            .lcout(\display2.prescaler_2_15 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_14 ),
            .carryout(\display2.prescaler_2_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_16_LC_14_13_7 .C_ON=1'b1;
    defparam \display2.prescaler_16_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_16_LC_14_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_16_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__13131),
            .in2(_gnd_net_),
            .in3(N__12888),
            .lcout(\display2.prescalerZ0Z_16 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_15 ),
            .carryout(\display2.prescaler_2_cry_16 ),
            .clk(N__14237),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_17_LC_14_14_0 .C_ON=1'b1;
    defparam \display2.prescaler_17_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_17_LC_14_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_17_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__13143),
            .in2(_gnd_net_),
            .in3(N__12885),
            .lcout(\display2.prescalerZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\display2.prescaler_2_cry_17 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_18_LC_14_14_1 .C_ON=1'b1;
    defparam \display2.prescaler_18_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_18_LC_14_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_18_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__13118),
            .in2(_gnd_net_),
            .in3(N__12882),
            .lcout(\display2.prescalerZ0Z_18 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_17 ),
            .carryout(\display2.prescaler_2_cry_18 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_19_LC_14_14_2 .C_ON=1'b1;
    defparam \display2.prescaler_19_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_19_LC_14_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \display2.prescaler_19_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12969),
            .in3(N__13032),
            .lcout(\display2.prescalerZ0Z_19 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_18 ),
            .carryout(\display2.prescaler_2_cry_19 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_20_LC_14_14_3 .C_ON=1'b1;
    defparam \display2.prescaler_20_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_20_LC_14_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_20_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__12993),
            .in2(_gnd_net_),
            .in3(N__13029),
            .lcout(\display2.prescalerZ0Z_20 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_19 ),
            .carryout(\display2.prescaler_2_cry_20 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_21_LC_14_14_4 .C_ON=1'b1;
    defparam \display2.prescaler_21_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_21_LC_14_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \display2.prescaler_21_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__13002),
            .in2(_gnd_net_),
            .in3(N__13026),
            .lcout(\display2.prescalerZ0Z_21 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_20 ),
            .carryout(\display2.prescaler_2_cry_21 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_22_LC_14_14_5 .C_ON=1'b1;
    defparam \display2.prescaler_22_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_22_LC_14_14_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \display2.prescaler_22_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12984),
            .in3(N__13023),
            .lcout(\display2.prescalerZ0Z_22 ),
            .ltout(),
            .carryin(\display2.prescaler_2_cry_21 ),
            .carryout(\display2.prescaler_2_cry_22 ),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_23_LC_14_14_6 .C_ON=1'b0;
    defparam \display2.prescaler_23_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_23_LC_14_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \display2.prescaler_23_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__13016),
            .in2(_gnd_net_),
            .in3(N__13020),
            .lcout(\display2.prescalerZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14230),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNIF8K21_19_LC_14_14_7 .C_ON=1'b0;
    defparam \display2.prescaler_RNIF8K21_19_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNIF8K21_19_LC_14_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display2.prescaler_RNIF8K21_19_LC_14_14_7  (
            .in0(N__13001),
            .in1(N__12992),
            .in2(N__12983),
            .in3(N__12965),
            .lcout(\display2.prescaler8_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNIDHIG_2_LC_15_12_3 .C_ON=1'b0;
    defparam \display2.prescaler_RNIDHIG_2_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNIDHIG_2_LC_15_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display2.prescaler_RNIDHIG_2_LC_15_12_3  (
            .in0(N__12956),
            .in1(N__12944),
            .in2(N__12933),
            .in3(N__12917),
            .lcout(\display2.prescaler8_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.digit_posn_LC_15_12_4 .C_ON=1'b0;
    defparam \display2.digit_posn_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \display2.digit_posn_LC_15_12_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \display2.digit_posn_LC_15_12_4  (
            .in0(N__13068),
            .in1(N__14032),
            .in2(N__13410),
            .in3(N__13994),
            .lcout(\display2.digit_posnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14250),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_0_LC_15_12_5 .C_ON=1'b0;
    defparam \display2.prescaler_0_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_0_LC_15_12_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \display2.prescaler_0_LC_15_12_5  (
            .in0(N__13995),
            .in1(N__13069),
            .in2(N__14042),
            .in3(N__13103),
            .lcout(\display2.prescalerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14250),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_1_LC_15_12_6 .C_ON=1'b0;
    defparam \display2.prescaler_1_LC_15_12_6 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_1_LC_15_12_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \display2.prescaler_1_LC_15_12_6  (
            .in0(N__13104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13205),
            .lcout(\display2.prescalerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14250),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNI6SG21_10_LC_15_13_0 .C_ON=1'b0;
    defparam \display2.prescaler_RNI6SG21_10_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNI6SG21_10_LC_15_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display2.prescaler_RNI6SG21_10_LC_15_13_0  (
            .in0(N__13284),
            .in1(N__13268),
            .in2(N__13257),
            .in3(N__13238),
            .lcout(),
            .ltout(\display2.prescaler8_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNI7PO13_1_LC_15_13_1 .C_ON=1'b0;
    defparam \display2.prescaler_RNI7PO13_1_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNI7PO13_1_LC_15_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \display2.prescaler_RNI7PO13_1_LC_15_13_1  (
            .in0(N__13227),
            .in1(N__13185),
            .in2(N__13218),
            .in3(N__13215),
            .lcout(\display2.prescaler8_21 ),
            .ltout(\display2.prescaler8_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNIQNE25_16_LC_15_13_2 .C_ON=1'b0;
    defparam \display2.prescaler_RNIQNE25_16_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNIQNE25_16_LC_15_13_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \display2.prescaler_RNIQNE25_16_LC_15_13_2  (
            .in0(N__13990),
            .in1(_gnd_net_),
            .in2(N__13209),
            .in3(N__13057),
            .lcout(\display2.prescaler8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNIHUHP_1_LC_15_13_3 .C_ON=1'b0;
    defparam \display2.prescaler_RNIHUHP_1_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNIHUHP_1_LC_15_13_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \display2.prescaler_RNIHUHP_1_LC_15_13_3  (
            .in0(N__13154),
            .in1(N__13172),
            .in2(N__13953),
            .in3(N__13204),
            .lcout(\display2.prescaler8_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_9_LC_15_13_4 .C_ON=1'b0;
    defparam \display2.prescaler_9_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_9_LC_15_13_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display2.prescaler_9_LC_15_13_4  (
            .in0(N__13993),
            .in1(N__14031),
            .in2(N__13081),
            .in3(N__13179),
            .lcout(\display2.prescalerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14243),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_14_LC_15_13_5 .C_ON=1'b0;
    defparam \display2.prescaler_14_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_14_LC_15_13_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \display2.prescaler_14_LC_15_13_5  (
            .in0(N__14030),
            .in1(N__13991),
            .in2(N__13073),
            .in3(N__13161),
            .lcout(\display2.prescalerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14243),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_RNI4M1U_16_LC_15_13_6 .C_ON=1'b0;
    defparam \display2.prescaler_RNI4M1U_16_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \display2.prescaler_RNI4M1U_16_LC_15_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \display2.prescaler_RNI4M1U_16_LC_15_13_6  (
            .in0(N__13142),
            .in1(N__13130),
            .in2(N__13119),
            .in3(N__13102),
            .lcout(\display2.prescaler8_17 ),
            .ltout(\display2.prescaler8_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.prescaler_15_LC_15_13_7 .C_ON=1'b0;
    defparam \display2.prescaler_15_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \display2.prescaler_15_LC_15_13_7 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \display2.prescaler_15_LC_15_13_7  (
            .in0(N__14049),
            .in1(N__14036),
            .in2(N__13998),
            .in3(N__13992),
            .lcout(\display2.prescalerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14243),
            .ce(),
            .sr(_gnd_net_));
    defparam \d1.sync_0_LC_16_8_7 .C_ON=1'b0;
    defparam \d1.sync_0_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \d1.sync_0_LC_16_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \d1.sync_0_LC_16_8_7  (
            .in0(N__13938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\d1.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14267),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.digit_data_3_LC_16_13_5 .C_ON=1'b0;
    defparam \display2.digit_data_3_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \display2.digit_data_3_LC_16_13_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \display2.digit_data_3_LC_16_13_5  (
            .in0(N__13344),
            .in1(N__13401),
            .in2(N__14465),
            .in3(N__13896),
            .lcout(\display2.digit_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14251),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.digit_data_2_LC_16_13_6 .C_ON=1'b0;
    defparam \display2.digit_data_2_LC_16_13_6 .SEQ_MODE=4'b1000;
    defparam \display2.digit_data_2_LC_16_13_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \display2.digit_data_2_LC_16_13_6  (
            .in0(N__13400),
            .in1(N__13343),
            .in2(N__14521),
            .in3(N__13794),
            .lcout(\display2.digit_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14251),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.digit_data_1_LC_16_14_6 .C_ON=1'b0;
    defparam \display2.digit_data_1_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \display2.digit_data_1_LC_16_14_6 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \display2.digit_data_1_LC_16_14_6  (
            .in0(N__13346),
            .in1(N__13412),
            .in2(N__14388),
            .in3(N__13683),
            .lcout(\display2.digit_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14244),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.digit_data_0_LC_16_14_7 .C_ON=1'b0;
    defparam \display2.digit_data_0_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \display2.digit_data_0_LC_16_14_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \display2.digit_data_0_LC_16_14_7  (
            .in0(N__13411),
            .in1(N__13345),
            .in2(N__14331),
            .in3(N__13554),
            .lcout(\display2.digit_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14244),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.DIGIT_e_0_LC_17_13_6 .C_ON=1'b0;
    defparam \display2.DIGIT_e_0_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \display2.DIGIT_e_0_LC_17_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \display2.DIGIT_e_0_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13416),
            .lcout(DIGIT_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14257),
            .ce(N__13353),
            .sr(_gnd_net_));
    defparam \d4.sync_0_LC_19_1_5 .C_ON=1'b0;
    defparam \d4.sync_0_LC_19_1_5 .SEQ_MODE=4'b1000;
    defparam \d4.sync_0_LC_19_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \d4.sync_0_LC_19_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13323),
            .lcout(\d4.syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14277),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_0_LC_23_13_7 .C_ON=1'b0;
    defparam \display2.decoder.SEG_0_LC_23_13_7 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_0_LC_23_13_7 .LUT_INIT=16'b0001011000110110;
    LogicCell40 \display2.decoder.SEG_0_LC_23_13_7  (
            .in0(N__14522),
            .in1(N__14476),
            .in2(N__14423),
            .in3(N__14350),
            .lcout(SEG2_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14274),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_5_LC_23_14_1 .C_ON=1'b0;
    defparam \display2.decoder.SEG_5_LC_23_14_1 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_5_LC_23_14_1 .LUT_INIT=16'b0011010100010111;
    LogicCell40 \display2.decoder.SEG_5_LC_23_14_1  (
            .in0(N__14541),
            .in1(N__14478),
            .in2(N__14405),
            .in3(N__14332),
            .lcout(SEG2_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14272),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_2_LC_24_13_1 .C_ON=1'b0;
    defparam \display2.decoder.SEG_2_LC_24_13_1 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_2_LC_24_13_1 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \display2.decoder.SEG_2_LC_24_13_1  (
            .in0(N__14352),
            .in1(N__14524),
            .in2(N__14477),
            .in3(N__14422),
            .lcout(SEG2_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14276),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_1_LC_24_13_4 .C_ON=1'b0;
    defparam \display2.decoder.SEG_1_LC_24_13_4 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_1_LC_24_13_4 .LUT_INIT=16'b0000011000100111;
    LogicCell40 \display2.decoder.SEG_1_LC_24_13_4  (
            .in0(N__14523),
            .in1(N__14461),
            .in2(N__14424),
            .in3(N__14351),
            .lcout(SEG2_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14276),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_4_LC_24_14_1 .C_ON=1'b0;
    defparam \display2.decoder.SEG_4_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_4_LC_24_14_1 .LUT_INIT=16'b0000111100111011;
    LogicCell40 \display2.decoder.SEG_4_LC_24_14_1  (
            .in0(N__14334),
            .in1(N__14395),
            .in2(N__14484),
            .in3(N__14543),
            .lcout(SEG2_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14275),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_3_LC_24_14_4 .C_ON=1'b0;
    defparam \display2.decoder.SEG_3_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_3_LC_24_14_4 .LUT_INIT=16'b0001011000110101;
    LogicCell40 \display2.decoder.SEG_3_LC_24_14_4  (
            .in0(N__14542),
            .in1(N__14479),
            .in2(N__14406),
            .in3(N__14333),
            .lcout(SEG2_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14275),
            .ce(),
            .sr(_gnd_net_));
    defparam \display2.decoder.SEG_6_LC_24_14_6 .C_ON=1'b0;
    defparam \display2.decoder.SEG_6_LC_24_14_6 .SEQ_MODE=4'b1000;
    defparam \display2.decoder.SEG_6_LC_24_14_6 .LUT_INIT=16'b0011011000110101;
    LogicCell40 \display2.decoder.SEG_6_LC_24_14_6  (
            .in0(N__14544),
            .in1(N__14480),
            .in2(N__14407),
            .in3(N__14335),
            .lcout(SEG2_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14275),
            .ce(),
            .sr(_gnd_net_));
endmodule // timer
